magic
tech sky130A
magscale 1 2
timestamp 1738079716
<< viali >>
rect 65717 63461 65751 63495
rect 66361 63325 66395 63359
rect 65625 61897 65659 61931
rect 66269 61693 66303 61727
rect 65625 60265 65659 60299
rect 66269 60061 66303 60095
rect 65625 58633 65659 58667
rect 66269 58429 66303 58463
rect 65625 57001 65659 57035
rect 66269 56797 66303 56831
rect 65625 55369 65659 55403
rect 66269 55233 66303 55267
rect 65809 53601 65843 53635
rect 67005 53533 67039 53567
rect 65625 53193 65659 53227
rect 66269 52989 66303 53023
rect 65625 52445 65659 52479
rect 65901 52445 65935 52479
rect 65625 51969 65659 52003
rect 66269 51901 66303 51935
rect 65625 50473 65659 50507
rect 66269 50337 66303 50371
rect 66361 50269 66395 50303
rect 65625 49589 65659 49623
rect 65625 49181 65659 49215
rect 65625 48841 65659 48875
rect 66269 48637 66303 48671
rect 65625 47209 65659 47243
rect 66361 47073 66395 47107
rect 66269 47005 66303 47039
rect 66637 46937 66671 46971
rect 65625 45509 65659 45543
rect 66269 45373 66303 45407
rect 65625 43945 65659 43979
rect 66269 43809 66303 43843
rect 66361 43741 66395 43775
rect 68017 42721 68051 42755
rect 65625 42653 65659 42687
rect 68661 42653 68695 42687
rect 65625 42313 65659 42347
rect 66269 42109 66303 42143
rect 66729 41769 66763 41803
rect 67373 41565 67407 41599
rect 65809 40885 65843 40919
rect 67097 40681 67131 40715
rect 65809 40545 65843 40579
rect 66821 40477 66855 40511
rect 67741 40477 67775 40511
rect 65625 40137 65659 40171
rect 66269 39933 66303 39967
rect 65625 39593 65659 39627
rect 66269 39389 66303 39423
rect 65625 39049 65659 39083
rect 66269 38845 66303 38879
rect 65625 38505 65659 38539
rect 66269 38301 66303 38335
rect 66269 37961 66303 37995
rect 65717 37757 65751 37791
rect 65625 37213 65659 37247
rect 66269 37213 66303 37247
rect 65625 36873 65659 36907
rect 66269 36669 66303 36703
rect 65625 36329 65659 36363
rect 66361 36329 66395 36363
rect 66269 36193 66303 36227
rect 67005 36125 67039 36159
rect 67097 35785 67131 35819
rect 66821 35717 66855 35751
rect 65625 35649 65659 35683
rect 67741 35581 67775 35615
rect 68017 35241 68051 35275
rect 67373 35105 67407 35139
rect 68569 35037 68603 35071
rect 65625 34969 65659 35003
rect 65625 34697 65659 34731
rect 67097 34697 67131 34731
rect 66361 34629 66395 34663
rect 66269 34493 66303 34527
rect 66913 34493 66947 34527
rect 67741 34493 67775 34527
rect 65625 34153 65659 34187
rect 66361 34153 66395 34187
rect 67097 34153 67131 34187
rect 66269 34017 66303 34051
rect 67005 33949 67039 33983
rect 67741 33949 67775 33983
rect 65625 33609 65659 33643
rect 66177 33405 66211 33439
rect 65625 33065 65659 33099
rect 66269 32861 66303 32895
rect 65625 32521 65659 32555
rect 66269 32317 66303 32351
rect 66269 31977 66303 32011
rect 65717 31773 65751 31807
rect 65625 31433 65659 31467
rect 66269 31229 66303 31263
rect 66269 30889 66303 30923
rect 65717 30685 65751 30719
rect 65625 30277 65659 30311
rect 66269 30141 66303 30175
rect 66269 29801 66303 29835
rect 65717 29597 65751 29631
rect 66269 29257 66303 29291
rect 65717 29121 65751 29155
rect 66913 28713 66947 28747
rect 65625 28441 65659 28475
rect 65625 28169 65659 28203
rect 66269 27965 66303 27999
rect 66637 27829 66671 27863
rect 66361 27557 66395 27591
rect 66913 27489 66947 27523
rect 66269 27421 66303 27455
rect 65625 27353 65659 27387
rect 67097 27081 67131 27115
rect 66545 27013 66579 27047
rect 65625 26945 65659 26979
rect 67741 26877 67775 26911
rect 65625 26537 65659 26571
rect 66269 26333 66303 26367
rect 65625 25993 65659 26027
rect 66269 25789 66303 25823
rect 65625 25449 65659 25483
rect 66269 25245 66303 25279
rect 66361 24769 66395 24803
rect 66269 24701 66303 24735
rect 67005 24701 67039 24735
rect 65625 24633 65659 24667
rect 65625 24361 65659 24395
rect 67005 24361 67039 24395
rect 66269 24225 66303 24259
rect 66361 24157 66395 24191
rect 65625 23817 65659 23851
rect 66361 23817 66395 23851
rect 67097 23817 67131 23851
rect 66269 23613 66303 23647
rect 66913 23613 66947 23647
rect 67741 23613 67775 23647
rect 67097 23273 67131 23307
rect 66361 23205 66395 23239
rect 66269 23137 66303 23171
rect 66913 23069 66947 23103
rect 67741 23069 67775 23103
rect 65625 23001 65659 23035
rect 65625 22729 65659 22763
rect 66269 22525 66303 22559
rect 66453 22049 66487 22083
rect 68661 22049 68695 22083
rect 70133 22049 70167 22083
rect 65809 21981 65843 22015
rect 69305 21981 69339 22015
rect 70777 21981 70811 22015
rect 65625 21641 65659 21675
rect 66269 21437 66303 21471
rect 68201 21097 68235 21131
rect 68845 20893 68879 20927
rect 67097 20553 67131 20587
rect 66361 20485 66395 20519
rect 67005 20417 67039 20451
rect 66269 20349 66303 20383
rect 67741 20349 67775 20383
rect 65625 20213 65659 20247
rect 65625 20009 65659 20043
rect 66269 19805 66303 19839
rect 66269 19465 66303 19499
rect 65717 19261 65751 19295
rect 66269 18921 66303 18955
rect 65717 18717 65751 18751
rect 65625 18377 65659 18411
rect 66269 18173 66303 18207
rect 66269 17833 66303 17867
rect 65717 17629 65751 17663
rect 65625 17289 65659 17323
rect 66361 17289 66395 17323
rect 66269 17085 66303 17119
rect 67005 17085 67039 17119
rect 66269 16609 66303 16643
rect 65625 16541 65659 16575
rect 65625 16201 65659 16235
rect 66269 15997 66303 16031
rect 65625 15657 65659 15691
rect 66269 15453 66303 15487
rect 65625 15113 65659 15147
rect 66269 14909 66303 14943
rect 65625 14569 65659 14603
rect 66269 14365 66303 14399
rect 65625 13481 65659 13515
rect 66269 13277 66303 13311
rect 65625 11849 65659 11883
rect 66269 11645 66303 11679
rect 39497 5865 39531 5899
rect 41705 5865 41739 5899
rect 49617 5865 49651 5899
rect 50721 5865 50755 5899
rect 53665 5865 53699 5899
rect 40417 5797 40451 5831
rect 29285 5729 29319 5763
rect 36369 5729 36403 5763
rect 46765 5729 46799 5763
rect 52193 5729 52227 5763
rect 60473 5729 60507 5763
rect 61025 5729 61059 5763
rect 28917 5661 28951 5695
rect 29101 5661 29135 5695
rect 29929 5661 29963 5695
rect 30665 5661 30699 5695
rect 31401 5661 31435 5695
rect 35725 5661 35759 5695
rect 36461 5661 36495 5695
rect 36737 5661 36771 5695
rect 37197 5661 37231 5695
rect 38117 5661 38151 5695
rect 38761 5661 38795 5695
rect 38853 5661 38887 5695
rect 39773 5661 39807 5695
rect 41061 5661 41095 5695
rect 45569 5661 45603 5695
rect 47501 5661 47535 5695
rect 48973 5661 49007 5695
rect 50077 5661 50111 5695
rect 50813 5661 50847 5695
rect 51549 5661 51583 5695
rect 53021 5661 53055 5695
rect 54401 5661 54435 5695
rect 55045 5661 55079 5695
rect 55229 5661 55263 5695
rect 56333 5661 56367 5695
rect 56701 5661 56735 5695
rect 57345 5661 57379 5695
rect 59369 5661 59403 5695
rect 29653 5593 29687 5627
rect 48697 5593 48731 5627
rect 30021 5525 30055 5559
rect 30849 5525 30883 5559
rect 37841 5525 37875 5559
rect 51457 5525 51491 5559
rect 60013 5525 60047 5559
rect 35725 5321 35759 5355
rect 37841 5321 37875 5355
rect 42165 5321 42199 5355
rect 42809 5321 42843 5355
rect 47317 5321 47351 5355
rect 48237 5321 48271 5355
rect 49065 5321 49099 5355
rect 49801 5321 49835 5355
rect 50537 5321 50571 5355
rect 54033 5321 54067 5355
rect 54769 5321 54803 5355
rect 56977 5321 57011 5355
rect 28917 5253 28951 5287
rect 46121 5253 46155 5287
rect 52009 5253 52043 5287
rect 29193 5185 29227 5219
rect 29377 5185 29411 5219
rect 32137 5185 32171 5219
rect 38577 5185 38611 5219
rect 41521 5185 41555 5219
rect 44097 5185 44131 5219
rect 44741 5185 44775 5219
rect 45477 5185 45511 5219
rect 55689 5185 55723 5219
rect 56425 5185 56459 5219
rect 26065 5117 26099 5151
rect 27445 5117 27479 5151
rect 28457 5117 28491 5151
rect 29929 5117 29963 5151
rect 30021 5117 30055 5151
rect 31125 5117 31159 5151
rect 33425 5117 33459 5151
rect 35081 5117 35115 5151
rect 37197 5117 37231 5151
rect 39221 5117 39255 5151
rect 40141 5117 40175 5151
rect 46673 5117 46707 5151
rect 47593 5117 47627 5151
rect 48421 5117 48455 5151
rect 49157 5117 49191 5151
rect 49893 5117 49927 5151
rect 50629 5117 50663 5151
rect 51273 5117 51307 5151
rect 51365 5117 51399 5151
rect 52653 5117 52687 5151
rect 53297 5117 53331 5151
rect 53389 5117 53423 5151
rect 54125 5117 54159 5151
rect 54861 5117 54895 5151
rect 26893 5049 26927 5083
rect 32413 5049 32447 5083
rect 40785 5049 40819 5083
rect 26709 4981 26743 5015
rect 27905 4981 27939 5015
rect 30665 4981 30699 5015
rect 31677 4981 31711 5015
rect 32873 4981 32907 5015
rect 45385 4981 45419 5015
rect 55505 4981 55539 5015
rect 56241 4981 56275 5015
rect 26157 4777 26191 4811
rect 31309 4777 31343 4811
rect 33793 4777 33827 4811
rect 35541 4777 35575 4811
rect 42901 4777 42935 4811
rect 26893 4709 26927 4743
rect 40601 4709 40635 4743
rect 25605 4641 25639 4675
rect 28365 4641 28399 4675
rect 34437 4641 34471 4675
rect 36185 4641 36219 4675
rect 42257 4641 42291 4675
rect 25053 4573 25087 4607
rect 26249 4573 26283 4607
rect 27997 4573 28031 4607
rect 28549 4573 28583 4607
rect 28641 4573 28675 4607
rect 29837 4573 29871 4607
rect 31217 4573 31251 4607
rect 31861 4573 31895 4607
rect 32965 4573 32999 4607
rect 33149 4573 33183 4607
rect 33977 4573 34011 4607
rect 34621 4573 34655 4607
rect 34897 4573 34931 4607
rect 36369 4573 36403 4607
rect 39957 4573 39991 4607
rect 41337 4573 41371 4607
rect 42993 4573 43027 4607
rect 44097 4573 44131 4607
rect 44741 4573 44775 4607
rect 45017 4573 45051 4607
rect 46121 4573 46155 4607
rect 46765 4573 46799 4607
rect 47225 4573 47259 4607
rect 47777 4573 47811 4607
rect 47869 4573 47903 4607
rect 51181 4573 51215 4607
rect 35265 4505 35299 4539
rect 36829 4505 36863 4539
rect 38025 4505 38059 4539
rect 43637 4505 43671 4539
rect 24501 4437 24535 4471
rect 27353 4437 27387 4471
rect 29285 4437 29319 4471
rect 30481 4437 30515 4471
rect 30573 4437 30607 4471
rect 32413 4437 32447 4471
rect 36737 4437 36771 4471
rect 37933 4437 37967 4471
rect 41981 4437 42015 4471
rect 45661 4437 45695 4471
rect 48513 4437 48547 4471
rect 51825 4437 51859 4471
rect 26893 4097 26927 4131
rect 27537 4097 27571 4131
rect 28917 4097 28951 4131
rect 29469 4097 29503 4131
rect 29653 4097 29687 4131
rect 30297 4097 30331 4131
rect 30941 4097 30975 4131
rect 32137 4097 32171 4131
rect 32689 4097 32723 4131
rect 37841 4097 37875 4131
rect 38945 4097 38979 4131
rect 43545 4097 43579 4131
rect 44281 4097 44315 4131
rect 47685 4097 47719 4131
rect 48237 4097 48271 4131
rect 53389 4097 53423 4131
rect 24593 4029 24627 4063
rect 25881 4029 25915 4063
rect 26617 4029 26651 4063
rect 27169 4029 27203 4063
rect 28181 4029 28215 4063
rect 30389 4029 30423 4063
rect 31769 4029 31803 4063
rect 33425 4029 33459 4063
rect 34161 4029 34195 4063
rect 34897 4029 34931 4063
rect 35633 4029 35667 4063
rect 36001 4029 36035 4063
rect 37657 4029 37691 4063
rect 38301 4029 38335 4063
rect 42165 4029 42199 4063
rect 42441 4029 42475 4063
rect 45477 4029 45511 4063
rect 52745 4029 52779 4063
rect 44097 3961 44131 3995
rect 46121 3961 46155 3995
rect 25237 3893 25271 3927
rect 25329 3893 25363 3927
rect 26065 3893 26099 3927
rect 28089 3893 28123 3927
rect 28825 3893 28859 3927
rect 31217 3893 31251 3927
rect 32873 3893 32907 3927
rect 33609 3893 33643 3927
rect 34345 3893 34379 3927
rect 35081 3893 35115 3927
rect 36645 3893 36679 3927
rect 41521 3893 41555 3927
rect 42993 3893 43027 3927
rect 44925 3893 44959 3927
rect 29285 3689 29319 3723
rect 31493 3689 31527 3723
rect 35357 3689 35391 3723
rect 42717 3689 42751 3723
rect 43453 3689 43487 3723
rect 49433 3689 49467 3723
rect 40877 3621 40911 3655
rect 25605 3553 25639 3587
rect 29837 3553 29871 3587
rect 34345 3553 34379 3587
rect 38945 3553 38979 3587
rect 41981 3553 42015 3587
rect 44005 3553 44039 3587
rect 45661 3553 45695 3587
rect 46489 3553 46523 3587
rect 47777 3553 47811 3587
rect 50905 3553 50939 3587
rect 64337 3553 64371 3587
rect 23581 3485 23615 3519
rect 24869 3485 24903 3519
rect 25697 3485 25731 3519
rect 26433 3485 26467 3519
rect 27813 3485 27847 3519
rect 27997 3485 28031 3519
rect 28733 3485 28767 3519
rect 30021 3485 30055 3519
rect 30665 3485 30699 3519
rect 30941 3485 30975 3519
rect 32229 3485 32263 3519
rect 32321 3485 32355 3519
rect 33057 3485 33091 3519
rect 34713 3485 34747 3519
rect 36001 3485 36035 3519
rect 36185 3485 36219 3519
rect 36829 3485 36863 3519
rect 37473 3485 37507 3519
rect 38393 3485 38427 3519
rect 39129 3485 39163 3519
rect 40325 3485 40359 3519
rect 40601 3485 40635 3519
rect 41337 3485 41371 3519
rect 43269 3485 43303 3519
rect 44649 3485 44683 3519
rect 45017 3485 45051 3519
rect 47225 3485 47259 3519
rect 47961 3485 47995 3519
rect 48605 3485 48639 3519
rect 49157 3485 49191 3519
rect 49617 3485 49651 3519
rect 50721 3485 50755 3519
rect 51733 3485 51767 3519
rect 53021 3485 53055 3519
rect 55873 3485 55907 3519
rect 57621 3485 57655 3519
rect 60473 3485 60507 3519
rect 64521 3485 64555 3519
rect 24593 3417 24627 3451
rect 27169 3417 27203 3451
rect 31585 3417 31619 3451
rect 36921 3417 36955 3451
rect 41061 3417 41095 3451
rect 44373 3417 44407 3451
rect 46305 3417 46339 3451
rect 52285 3417 52319 3451
rect 58633 3417 58667 3451
rect 60841 3417 60875 3451
rect 24133 3349 24167 3383
rect 24961 3349 24995 3383
rect 26341 3349 26375 3383
rect 27077 3349 27111 3383
rect 28549 3349 28583 3383
rect 30113 3349 30147 3383
rect 32965 3349 32999 3383
rect 33701 3349 33735 3383
rect 33793 3349 33827 3383
rect 35449 3349 35483 3383
rect 37841 3349 37875 3383
rect 41889 3349 41923 3383
rect 42625 3349 42659 3383
rect 45569 3349 45603 3383
rect 47041 3349 47075 3383
rect 48513 3349 48547 3383
rect 50077 3349 50111 3383
rect 51457 3349 51491 3383
rect 52377 3349 52411 3383
rect 55229 3349 55263 3383
rect 58173 3349 58207 3383
rect 58541 3349 58575 3383
rect 23029 3145 23063 3179
rect 31861 3145 31895 3179
rect 32597 3145 32631 3179
rect 34713 3145 34747 3179
rect 35449 3145 35483 3179
rect 36277 3145 36311 3179
rect 38025 3145 38059 3179
rect 39773 3145 39807 3179
rect 42349 3145 42383 3179
rect 45293 3145 45327 3179
rect 46857 3145 46891 3179
rect 47501 3145 47535 3179
rect 48973 3145 49007 3179
rect 52193 3145 52227 3179
rect 52653 3145 52687 3179
rect 57345 3145 57379 3179
rect 60749 3145 60783 3179
rect 24501 3077 24535 3111
rect 29285 3077 29319 3111
rect 31125 3077 31159 3111
rect 32413 3077 32447 3111
rect 33333 3077 33367 3111
rect 52285 3077 52319 3111
rect 57437 3077 57471 3111
rect 62221 3077 62255 3111
rect 68293 3077 68327 3111
rect 23765 3009 23799 3043
rect 25237 3009 25271 3043
rect 26709 3009 26743 3043
rect 29745 3009 29779 3043
rect 31217 3009 31251 3043
rect 33241 3009 33275 3043
rect 33885 3009 33919 3043
rect 34897 3009 34931 3043
rect 35633 3009 35667 3043
rect 36829 3009 36863 3043
rect 39865 3009 39899 3043
rect 40877 3009 40911 3043
rect 42073 3009 42107 3043
rect 43821 3009 43855 3043
rect 47041 3009 47075 3043
rect 48237 3009 48271 3043
rect 49709 3009 49743 3043
rect 50445 3009 50479 3043
rect 53205 3009 53239 3043
rect 53481 3009 53515 3043
rect 55597 3009 55631 3043
rect 58541 3009 58575 3043
rect 59185 3009 59219 3043
rect 62589 3009 62623 3043
rect 64521 3009 64555 3043
rect 68569 3009 68603 3043
rect 69581 3009 69615 3043
rect 22385 2941 22419 2975
rect 23121 2941 23155 2975
rect 23857 2941 23891 2975
rect 25329 2941 25363 2975
rect 27169 2941 27203 2975
rect 27721 2941 27755 2975
rect 29561 2941 29595 2975
rect 30481 2941 30515 2975
rect 32137 2941 32171 2975
rect 34161 2941 34195 2975
rect 37289 2941 37323 2975
rect 37933 2941 37967 2975
rect 38577 2941 38611 2975
rect 39405 2941 39439 2975
rect 40233 2941 40267 2975
rect 42993 2941 43027 2975
rect 43729 2941 43763 2975
rect 44649 2941 44683 2975
rect 45201 2941 45235 2975
rect 45845 2941 45879 2975
rect 46121 2941 46155 2975
rect 46673 2941 46707 2975
rect 48053 2941 48087 2975
rect 48789 2941 48823 2975
rect 49525 2941 49559 2975
rect 51825 2941 51859 2975
rect 54033 2941 54067 2975
rect 54125 2941 54159 2975
rect 54861 2941 54895 2975
rect 56333 2941 56367 2975
rect 57805 2941 57839 2975
rect 59277 2941 59311 2975
rect 60013 2941 60047 2975
rect 61393 2941 61427 2975
rect 61577 2941 61611 2975
rect 63233 2941 63267 2975
rect 63785 2941 63819 2975
rect 63877 2941 63911 2975
rect 65257 2941 65291 2975
rect 65717 2941 65751 2975
rect 66269 2941 66303 2975
rect 66361 2941 66395 2975
rect 67189 2941 67223 2975
rect 69029 2941 69063 2975
rect 69673 2941 69707 2975
rect 71053 2941 71087 2975
rect 71329 2941 71363 2975
rect 25973 2873 26007 2907
rect 43085 2873 43119 2907
rect 50353 2873 50387 2907
rect 55505 2873 55539 2907
rect 62129 2873 62163 2907
rect 70317 2873 70351 2907
rect 24593 2805 24627 2839
rect 26065 2805 26099 2839
rect 27813 2805 27847 2839
rect 30389 2805 30423 2839
rect 36185 2805 36219 2839
rect 38761 2805 38795 2839
rect 40785 2805 40819 2839
rect 41521 2805 41555 2839
rect 41981 2805 42015 2839
rect 44465 2805 44499 2839
rect 51089 2805 51123 2839
rect 51181 2805 51215 2839
rect 54769 2805 54803 2839
rect 56241 2805 56275 2839
rect 56977 2805 57011 2839
rect 58449 2805 58483 2839
rect 59921 2805 59955 2839
rect 60657 2805 60691 2839
rect 64613 2805 64647 2839
rect 67005 2805 67039 2839
rect 67741 2805 67775 2839
rect 70409 2805 70443 2839
rect 71881 2805 71915 2839
rect 22661 2601 22695 2635
rect 23397 2601 23431 2635
rect 26709 2601 26743 2635
rect 28273 2601 28307 2635
rect 29469 2601 29503 2635
rect 29653 2601 29687 2635
rect 30113 2601 30147 2635
rect 32229 2601 32263 2635
rect 34437 2601 34471 2635
rect 35449 2601 35483 2635
rect 36921 2601 36955 2635
rect 37657 2601 37691 2635
rect 41245 2601 41279 2635
rect 43361 2601 43395 2635
rect 44925 2601 44959 2635
rect 45661 2601 45695 2635
rect 46397 2601 46431 2635
rect 48605 2601 48639 2635
rect 49433 2601 49467 2635
rect 50813 2601 50847 2635
rect 51549 2601 51583 2635
rect 53021 2601 53055 2635
rect 54769 2601 54803 2635
rect 65533 2601 65567 2635
rect 66269 2601 66303 2635
rect 69121 2601 69155 2635
rect 71421 2601 71455 2635
rect 30021 2533 30055 2567
rect 31493 2533 31527 2567
rect 33701 2533 33735 2567
rect 55965 2533 55999 2567
rect 59829 2533 59863 2567
rect 61853 2533 61887 2567
rect 63325 2533 63359 2567
rect 64429 2533 64463 2567
rect 22845 2465 22879 2499
rect 24685 2465 24719 2499
rect 25237 2465 25271 2499
rect 26065 2465 26099 2499
rect 28733 2465 28767 2499
rect 30757 2465 30791 2499
rect 30941 2465 30975 2499
rect 31677 2465 31711 2499
rect 33793 2465 33827 2499
rect 34897 2465 34931 2499
rect 36277 2465 36311 2499
rect 38393 2465 38427 2499
rect 38761 2465 38795 2499
rect 41797 2465 41831 2499
rect 42717 2465 42751 2499
rect 43453 2465 43487 2499
rect 46949 2465 46983 2499
rect 47133 2465 47167 2499
rect 50629 2465 50663 2499
rect 52101 2465 52135 2499
rect 54309 2465 54343 2499
rect 55229 2465 55263 2499
rect 56609 2465 56643 2499
rect 57253 2465 57287 2499
rect 58909 2465 58943 2499
rect 60381 2465 60415 2499
rect 61117 2465 61151 2499
rect 62589 2465 62623 2499
rect 64981 2465 65015 2499
rect 66821 2465 66855 2499
rect 67005 2465 67039 2499
rect 68477 2465 68511 2499
rect 70133 2465 70167 2499
rect 70685 2465 70719 2499
rect 72249 2465 72283 2499
rect 22109 2397 22143 2431
rect 24133 2397 24167 2431
rect 24317 2397 24351 2431
rect 25421 2397 25455 2431
rect 28181 2397 28215 2431
rect 28457 2397 28491 2431
rect 29285 2397 29319 2431
rect 32321 2397 32355 2431
rect 33057 2397 33091 2431
rect 35541 2397 35575 2431
rect 37105 2397 37139 2431
rect 37749 2397 37783 2431
rect 40417 2397 40451 2431
rect 40509 2397 40543 2431
rect 41061 2397 41095 2431
rect 41981 2397 42015 2431
rect 44097 2397 44131 2431
rect 44189 2397 44223 2431
rect 45569 2397 45603 2431
rect 46213 2397 46247 2431
rect 47777 2397 47811 2431
rect 47869 2397 47903 2431
rect 49249 2397 49283 2431
rect 49617 2397 49651 2431
rect 50077 2397 50111 2431
rect 51365 2397 51399 2431
rect 52285 2397 52319 2431
rect 53665 2397 53699 2431
rect 53757 2397 53791 2431
rect 54861 2397 54895 2431
rect 57529 2397 57563 2431
rect 58173 2397 58207 2431
rect 58725 2397 58759 2431
rect 62405 2397 62439 2431
rect 63877 2397 63911 2431
rect 66085 2397 66119 2431
rect 67741 2397 67775 2431
rect 69213 2397 69247 2431
rect 70409 2397 70443 2431
rect 71329 2397 71363 2431
rect 71973 2397 72007 2431
rect 26985 2329 27019 2363
rect 29653 2329 29687 2363
rect 44465 2329 44499 2363
rect 55873 2329 55907 2363
rect 60013 2329 60047 2363
rect 23489 2261 23523 2295
rect 24501 2261 24535 2295
rect 25973 2261 26007 2295
rect 32965 2261 32999 2295
rect 36185 2261 36219 2295
rect 39405 2261 39439 2295
rect 39773 2261 39807 2295
rect 42625 2261 42659 2295
rect 48513 2261 48547 2295
rect 52929 2261 52963 2295
rect 56701 2261 56735 2295
rect 58081 2261 58115 2295
rect 59553 2261 59587 2295
rect 61025 2261 61059 2295
rect 61761 2261 61795 2295
rect 63233 2261 63267 2295
rect 67649 2261 67683 2295
rect 68385 2261 68419 2295
rect 69857 2261 69891 2295
rect 72801 2261 72835 2295
rect 21557 2057 21591 2091
rect 25973 2057 26007 2091
rect 26985 2057 27019 2091
rect 36277 2057 36311 2091
rect 37013 2057 37047 2091
rect 39037 2057 39071 2091
rect 39773 2057 39807 2091
rect 41245 2057 41279 2091
rect 45385 2057 45419 2091
rect 46121 2057 46155 2091
rect 55965 2057 55999 2091
rect 58449 2057 58483 2091
rect 60473 2057 60507 2091
rect 61945 2057 61979 2091
rect 66085 2057 66119 2091
rect 70133 2057 70167 2091
rect 22753 1989 22787 2023
rect 49433 1989 49467 2023
rect 50537 1989 50571 2023
rect 52653 1989 52687 2023
rect 68385 1989 68419 2023
rect 71145 1989 71179 2023
rect 73445 1989 73479 2023
rect 22201 1921 22235 1955
rect 23489 1921 23523 1955
rect 24317 1921 24351 1955
rect 25789 1921 25823 1955
rect 26893 1921 26927 1955
rect 27261 1921 27295 1955
rect 29009 1921 29043 1955
rect 30205 1921 30239 1955
rect 31861 1921 31895 1955
rect 33701 1921 33735 1955
rect 35541 1921 35575 1955
rect 35725 1921 35759 1955
rect 36461 1921 36495 1955
rect 38577 1921 38611 1955
rect 39589 1921 39623 1955
rect 40325 1921 40359 1955
rect 41797 1921 41831 1955
rect 43821 1921 43855 1955
rect 45293 1921 45327 1955
rect 45937 1921 45971 1955
rect 46857 1921 46891 1955
rect 47501 1921 47535 1955
rect 49341 1921 49375 1955
rect 49985 1921 50019 1955
rect 50169 1921 50203 1955
rect 52101 1921 52135 1955
rect 53205 1921 53239 1955
rect 54861 1921 54895 1955
rect 54953 1921 54987 1955
rect 55505 1921 55539 1955
rect 56057 1921 56091 1955
rect 57621 1921 57655 1955
rect 60381 1921 60415 1955
rect 61209 1921 61243 1955
rect 62497 1921 62531 1955
rect 63325 1921 63359 1955
rect 64613 1921 64647 1955
rect 66821 1921 66855 1955
rect 68109 1921 68143 1955
rect 68661 1921 68695 1955
rect 70685 1921 70719 1955
rect 70869 1921 70903 1955
rect 71605 1921 71639 1955
rect 73721 1921 73755 1955
rect 21005 1853 21039 1887
rect 23581 1853 23615 1887
rect 25513 1853 25547 1887
rect 26157 1853 26191 1887
rect 28457 1853 28491 1887
rect 30665 1853 30699 1887
rect 32505 1853 32539 1887
rect 34345 1853 34379 1887
rect 37381 1853 37415 1887
rect 41061 1853 41095 1887
rect 42625 1853 42659 1887
rect 44189 1853 44223 1887
rect 46673 1853 46707 1887
rect 48145 1853 48179 1887
rect 50905 1853 50939 1887
rect 53665 1853 53699 1887
rect 56425 1853 56459 1887
rect 57805 1853 57839 1887
rect 59185 1853 59219 1887
rect 61025 1853 61059 1887
rect 63601 1853 63635 1887
rect 65073 1853 65107 1887
rect 66637 1853 66671 1887
rect 69121 1853 69155 1887
rect 71881 1853 71915 1887
rect 24225 1785 24259 1819
rect 61853 1785 61887 1819
rect 22845 1717 22879 1751
rect 26709 1717 26743 1751
rect 40509 1717 40543 1751
rect 47041 1717 47075 1751
rect 47685 1717 47719 1751
rect 67465 1717 67499 1751
rect 23489 1513 23523 1547
rect 32689 1513 32723 1547
rect 35449 1513 35483 1547
rect 43821 1513 43855 1547
rect 46673 1513 46707 1547
rect 67741 1513 67775 1547
rect 73997 1513 74031 1547
rect 21925 1445 21959 1479
rect 61853 1445 61887 1479
rect 22845 1377 22879 1411
rect 49525 1377 49559 1411
rect 64981 1377 65015 1411
rect 68569 1377 68603 1411
rect 71145 1377 71179 1411
rect 74641 1377 74675 1411
rect 20269 1309 20303 1343
rect 21005 1309 21039 1343
rect 21741 1309 21775 1343
rect 22017 1309 22051 1343
rect 24133 1309 24167 1343
rect 25605 1309 25639 1343
rect 26433 1309 26467 1343
rect 26709 1309 26743 1343
rect 27169 1309 27203 1343
rect 27813 1309 27847 1343
rect 29285 1309 29319 1343
rect 29837 1309 29871 1343
rect 31769 1309 31803 1343
rect 32137 1309 32171 1343
rect 32965 1309 32999 1343
rect 34897 1309 34931 1343
rect 36921 1309 36955 1343
rect 37565 1309 37599 1343
rect 39405 1309 39439 1343
rect 41153 1309 41187 1343
rect 41797 1309 41831 1343
rect 43729 1309 43763 1343
rect 44465 1309 44499 1343
rect 46397 1309 46431 1343
rect 47225 1309 47259 1343
rect 48881 1309 48915 1343
rect 51457 1309 51491 1343
rect 51549 1309 51583 1343
rect 52101 1309 52135 1343
rect 54033 1309 54067 1343
rect 54677 1309 54711 1343
rect 56517 1309 56551 1343
rect 56701 1309 56735 1343
rect 57253 1309 57287 1343
rect 59093 1309 59127 1343
rect 59277 1309 59311 1343
rect 59829 1309 59863 1343
rect 61761 1309 61795 1343
rect 62405 1309 62439 1343
rect 63141 1309 63175 1343
rect 64429 1309 64463 1343
rect 65901 1309 65935 1343
rect 67465 1309 67499 1343
rect 68201 1309 68235 1343
rect 69581 1309 69615 1343
rect 70133 1309 70167 1343
rect 70777 1309 70811 1343
rect 72157 1309 72191 1343
rect 72709 1309 72743 1343
rect 73261 1309 73295 1343
rect 73813 1309 73847 1343
rect 24593 1241 24627 1275
rect 28365 1241 28399 1275
rect 30941 1241 30975 1275
rect 33977 1241 34011 1275
rect 35725 1241 35759 1275
rect 38393 1241 38427 1275
rect 40049 1241 40083 1275
rect 41245 1241 41279 1275
rect 42533 1241 42567 1275
rect 45385 1241 45419 1275
rect 47685 1241 47719 1275
rect 48973 1241 49007 1275
rect 50261 1241 50295 1275
rect 52837 1241 52871 1275
rect 55413 1241 55447 1275
rect 57989 1241 58023 1275
rect 60565 1241 60599 1275
rect 63877 1241 63911 1275
rect 66821 1241 66855 1275
rect 20821 1173 20855 1207
rect 21557 1173 21591 1207
rect 22661 1173 22695 1207
rect 23397 1173 23431 1207
rect 30389 1173 30423 1207
rect 38117 1173 38151 1207
rect 54125 1173 54159 1207
<< metal1 >>
rect 65320 85978 74980 86000
rect 65320 85926 74210 85978
rect 74262 85926 74274 85978
rect 74326 85926 74338 85978
rect 74390 85926 74402 85978
rect 74454 85926 74466 85978
rect 74518 85926 74980 85978
rect 65320 85904 74980 85926
rect 65320 85434 74980 85456
rect 65320 85382 71858 85434
rect 71910 85382 71922 85434
rect 71974 85382 71986 85434
rect 72038 85382 72050 85434
rect 72102 85382 72114 85434
rect 72166 85382 74980 85434
rect 65320 85360 74980 85382
rect 65320 84890 74980 84912
rect 65320 84838 74210 84890
rect 74262 84838 74274 84890
rect 74326 84838 74338 84890
rect 74390 84838 74402 84890
rect 74454 84838 74466 84890
rect 74518 84838 74980 84890
rect 65320 84816 74980 84838
rect 65320 84346 74980 84368
rect 65320 84294 71858 84346
rect 71910 84294 71922 84346
rect 71974 84294 71986 84346
rect 72038 84294 72050 84346
rect 72102 84294 72114 84346
rect 72166 84294 74980 84346
rect 65320 84272 74980 84294
rect 64874 84232 64880 84244
rect 63236 84204 64880 84232
rect 64874 84192 64880 84204
rect 64932 84192 64938 84244
rect 65320 83802 74980 83824
rect 65320 83750 74210 83802
rect 74262 83750 74274 83802
rect 74326 83750 74338 83802
rect 74390 83750 74402 83802
rect 74454 83750 74466 83802
rect 74518 83750 74980 83802
rect 65320 83728 74980 83750
rect 65320 83258 74980 83280
rect 63236 83144 63264 83256
rect 65320 83206 71858 83258
rect 71910 83206 71922 83258
rect 71974 83206 71986 83258
rect 72038 83206 72050 83258
rect 72102 83206 72114 83258
rect 72166 83206 74980 83258
rect 65320 83184 74980 83206
rect 65702 83144 65708 83156
rect 63236 83116 65708 83144
rect 65702 83104 65708 83116
rect 65760 83104 65766 83156
rect 71682 83008 71688 83020
rect 63236 82980 71688 83008
rect 71682 82968 71688 82980
rect 71740 82968 71746 83020
rect 65320 82714 74980 82736
rect 65320 82662 74210 82714
rect 74262 82662 74274 82714
rect 74326 82662 74338 82714
rect 74390 82662 74402 82714
rect 74454 82662 74466 82714
rect 74518 82662 74980 82714
rect 65320 82640 74980 82662
rect 65320 82170 74980 82192
rect 65320 82118 71858 82170
rect 71910 82118 71922 82170
rect 71974 82118 71986 82170
rect 72038 82118 72050 82170
rect 72102 82118 72114 82170
rect 72166 82118 74980 82170
rect 65320 82096 74980 82118
rect 63236 81784 63264 82052
rect 64874 81784 64880 81796
rect 63236 81756 64880 81784
rect 64874 81744 64880 81756
rect 64932 81744 64938 81796
rect 65320 81626 74980 81648
rect 65320 81574 74210 81626
rect 74262 81574 74274 81626
rect 74326 81574 74338 81626
rect 74390 81574 74402 81626
rect 74454 81574 74466 81626
rect 74518 81574 74980 81626
rect 65320 81552 74980 81574
rect 65320 81082 74980 81104
rect 63236 80968 63264 81076
rect 65320 81030 71858 81082
rect 71910 81030 71922 81082
rect 71974 81030 71986 81082
rect 72038 81030 72050 81082
rect 72102 81030 72114 81082
rect 72166 81030 74980 81082
rect 65320 81008 74980 81030
rect 65518 80968 65524 80980
rect 63236 80940 65524 80968
rect 65518 80928 65524 80940
rect 65576 80928 65582 80980
rect 70670 80832 70676 80844
rect 63236 80804 70676 80832
rect 70670 80792 70676 80804
rect 70728 80792 70734 80844
rect 65320 80538 74980 80560
rect 65320 80486 74210 80538
rect 74262 80486 74274 80538
rect 74326 80486 74338 80538
rect 74390 80486 74402 80538
rect 74454 80486 74466 80538
rect 74518 80486 74980 80538
rect 65320 80464 74980 80486
rect 65320 79994 74980 80016
rect 65320 79942 71858 79994
rect 71910 79942 71922 79994
rect 71974 79942 71986 79994
rect 72038 79942 72050 79994
rect 72102 79942 72114 79994
rect 72166 79942 74980 79994
rect 65320 79920 74980 79942
rect 64874 79880 64880 79892
rect 63236 79852 64880 79880
rect 64874 79840 64880 79852
rect 64932 79840 64938 79892
rect 65320 79450 74980 79472
rect 65320 79398 74210 79450
rect 74262 79398 74274 79450
rect 74326 79398 74338 79450
rect 74390 79398 74402 79450
rect 74454 79398 74466 79450
rect 74518 79398 74980 79450
rect 65320 79376 74980 79398
rect 65320 78906 74980 78928
rect 63236 78724 63264 78896
rect 65320 78854 71858 78906
rect 71910 78854 71922 78906
rect 71974 78854 71986 78906
rect 72038 78854 72050 78906
rect 72102 78854 72114 78906
rect 72166 78854 74980 78906
rect 65320 78832 74980 78854
rect 65610 78724 65616 78736
rect 63236 78696 65616 78724
rect 65610 78684 65616 78696
rect 65668 78684 65674 78736
rect 68646 78656 68652 78668
rect 63236 78628 68652 78656
rect 68646 78616 68652 78628
rect 68704 78616 68710 78668
rect 65320 78362 74980 78384
rect 65320 78310 74210 78362
rect 74262 78310 74274 78362
rect 74326 78310 74338 78362
rect 74390 78310 74402 78362
rect 74454 78310 74466 78362
rect 74518 78310 74980 78362
rect 65320 78288 74980 78310
rect 65320 77818 74980 77840
rect 65320 77766 71858 77818
rect 71910 77766 71922 77818
rect 71974 77766 71986 77818
rect 72038 77766 72050 77818
rect 72102 77766 72114 77818
rect 72166 77766 74980 77818
rect 65320 77744 74980 77766
rect 64874 77704 64880 77716
rect 63236 77676 64880 77704
rect 64874 77664 64880 77676
rect 64932 77664 64938 77716
rect 65320 77274 74980 77296
rect 65320 77222 74210 77274
rect 74262 77222 74274 77274
rect 74326 77222 74338 77274
rect 74390 77222 74402 77274
rect 74454 77222 74466 77274
rect 74518 77222 74980 77274
rect 65320 77200 74980 77222
rect 65320 76730 74980 76752
rect 63236 76548 63264 76716
rect 65320 76678 71858 76730
rect 71910 76678 71922 76730
rect 71974 76678 71986 76730
rect 72038 76678 72050 76730
rect 72102 76678 72114 76730
rect 72166 76678 74980 76730
rect 65320 76656 74980 76678
rect 65334 76548 65340 76560
rect 63236 76520 65340 76548
rect 65334 76508 65340 76520
rect 65392 76508 65398 76560
rect 68094 76480 68100 76492
rect 63236 76452 68100 76480
rect 68094 76440 68100 76452
rect 68152 76440 68158 76492
rect 65320 76186 74980 76208
rect 65320 76134 74210 76186
rect 74262 76134 74274 76186
rect 74326 76134 74338 76186
rect 74390 76134 74402 76186
rect 74454 76134 74466 76186
rect 74518 76134 74980 76186
rect 65320 76112 74980 76134
rect 65320 75642 74980 75664
rect 65320 75590 71858 75642
rect 71910 75590 71922 75642
rect 71974 75590 71986 75642
rect 72038 75590 72050 75642
rect 72102 75590 72114 75642
rect 72166 75590 74980 75642
rect 65320 75568 74980 75590
rect 63236 75188 63264 75512
rect 64874 75188 64880 75200
rect 63236 75160 64880 75188
rect 64874 75148 64880 75160
rect 64932 75148 64938 75200
rect 65320 75098 74980 75120
rect 65320 75046 74210 75098
rect 74262 75046 74274 75098
rect 74326 75046 74338 75098
rect 74390 75046 74402 75098
rect 74454 75046 74466 75098
rect 74518 75046 74980 75098
rect 65320 75024 74980 75046
rect 65426 74644 65432 74656
rect 63236 74616 65432 74644
rect 63236 74536 63264 74616
rect 65426 74604 65432 74616
rect 65484 74604 65490 74656
rect 65320 74554 74980 74576
rect 65320 74502 71858 74554
rect 71910 74502 71922 74554
rect 71974 74502 71986 74554
rect 72038 74502 72050 74554
rect 72102 74502 72114 74554
rect 72166 74502 74980 74554
rect 65320 74480 74980 74502
rect 63236 74100 63264 74284
rect 65886 74100 65892 74112
rect 63236 74072 65892 74100
rect 65886 74060 65892 74072
rect 65944 74060 65950 74112
rect 65320 74010 74980 74032
rect 65320 73958 74210 74010
rect 74262 73958 74274 74010
rect 74326 73958 74338 74010
rect 74390 73958 74402 74010
rect 74454 73958 74466 74010
rect 74518 73958 74980 74010
rect 65320 73936 74980 73958
rect 65320 73466 74980 73488
rect 65320 73414 71858 73466
rect 71910 73414 71922 73466
rect 71974 73414 71986 73466
rect 72038 73414 72050 73466
rect 72102 73414 72114 73466
rect 72166 73414 74980 73466
rect 65320 73392 74980 73414
rect 63236 73216 63264 73332
rect 64874 73216 64880 73228
rect 63236 73188 64880 73216
rect 64874 73176 64880 73188
rect 64932 73176 64938 73228
rect 65320 72922 74980 72944
rect 65320 72870 74210 72922
rect 74262 72870 74274 72922
rect 74326 72870 74338 72922
rect 74390 72870 74402 72922
rect 74454 72870 74466 72922
rect 74518 72870 74980 72922
rect 65320 72848 74980 72870
rect 65320 72378 74980 72400
rect 63236 72196 63264 72356
rect 65320 72326 71858 72378
rect 71910 72326 71922 72378
rect 71974 72326 71986 72378
rect 72038 72326 72050 72378
rect 72102 72326 72114 72378
rect 72166 72326 74980 72378
rect 65320 72304 74980 72326
rect 65150 72196 65156 72208
rect 63236 72168 65156 72196
rect 65150 72156 65156 72168
rect 65208 72156 65214 72208
rect 63236 71788 63264 72104
rect 65320 71834 74980 71856
rect 64598 71788 64604 71800
rect 63236 71760 64604 71788
rect 64598 71748 64604 71760
rect 64656 71748 64662 71800
rect 65320 71782 74210 71834
rect 74262 71782 74274 71834
rect 74326 71782 74338 71834
rect 74390 71782 74402 71834
rect 74454 71782 74466 71834
rect 74518 71782 74980 71834
rect 65320 71760 74980 71782
rect 65320 71290 74980 71312
rect 65320 71238 71858 71290
rect 71910 71238 71922 71290
rect 71974 71238 71986 71290
rect 72038 71238 72050 71290
rect 72102 71238 72114 71290
rect 72166 71238 74980 71290
rect 65320 71216 74980 71238
rect 63236 71148 63816 71176
rect 63788 71108 63816 71148
rect 64874 71108 64880 71120
rect 63788 71080 64880 71108
rect 64874 71068 64880 71080
rect 64932 71068 64938 71120
rect 65320 70746 74980 70768
rect 65320 70694 74210 70746
rect 74262 70694 74274 70746
rect 74326 70694 74338 70746
rect 74390 70694 74402 70746
rect 74454 70694 74466 70746
rect 74518 70694 74980 70746
rect 65320 70672 74980 70694
rect 65320 70202 74980 70224
rect 63236 70020 63264 70176
rect 65320 70150 71858 70202
rect 71910 70150 71922 70202
rect 71974 70150 71986 70202
rect 72038 70150 72050 70202
rect 72102 70150 72114 70202
rect 72166 70150 74980 70202
rect 65320 70128 74980 70150
rect 65242 70020 65248 70032
rect 63236 69992 65248 70020
rect 65242 69980 65248 69992
rect 65300 69980 65306 70032
rect 71130 69952 71136 69964
rect 63236 69924 71136 69952
rect 71130 69912 71136 69924
rect 71188 69912 71194 69964
rect 65320 69658 74980 69680
rect 65320 69606 74210 69658
rect 74262 69606 74274 69658
rect 74326 69606 74338 69658
rect 74390 69606 74402 69658
rect 74454 69606 74466 69658
rect 74518 69606 74980 69658
rect 65320 69584 74980 69606
rect 65320 69114 74980 69136
rect 65320 69062 71858 69114
rect 71910 69062 71922 69114
rect 71974 69062 71986 69114
rect 72038 69062 72050 69114
rect 72102 69062 72114 69114
rect 72166 69062 74980 69114
rect 65320 69040 74980 69062
rect 63144 68972 63816 69000
rect 63788 68932 63816 68972
rect 64874 68932 64880 68944
rect 63788 68904 64880 68932
rect 64874 68892 64880 68904
rect 64932 68932 64938 68944
rect 65794 68932 65800 68944
rect 64932 68904 65800 68932
rect 64932 68892 64938 68904
rect 65794 68892 65800 68904
rect 65852 68892 65858 68944
rect 65320 68570 74980 68592
rect 65320 68518 74210 68570
rect 74262 68518 74274 68570
rect 74326 68518 74338 68570
rect 74390 68518 74402 68570
rect 74454 68518 74466 68570
rect 74518 68518 74980 68570
rect 65320 68496 74980 68518
rect 65320 68026 74980 68048
rect 63236 67844 63264 67996
rect 65320 67974 71858 68026
rect 71910 67974 71922 68026
rect 71974 67974 71986 68026
rect 72038 67974 72050 68026
rect 72102 67974 72114 68026
rect 72166 67974 74980 68026
rect 65320 67952 74980 67974
rect 65058 67844 65064 67856
rect 63236 67816 65064 67844
rect 65058 67804 65064 67816
rect 65116 67804 65122 67856
rect 72786 67776 72792 67788
rect 63236 67748 72792 67776
rect 63236 67744 63264 67748
rect 72786 67736 72792 67748
rect 72844 67736 72850 67788
rect 65320 67482 74980 67504
rect 65320 67430 74210 67482
rect 74262 67430 74274 67482
rect 74326 67430 74338 67482
rect 74390 67430 74402 67482
rect 74454 67430 74466 67482
rect 74518 67430 74980 67482
rect 65320 67408 74980 67430
rect 65320 66938 74980 66960
rect 65320 66886 71858 66938
rect 71910 66886 71922 66938
rect 71974 66886 71986 66938
rect 72038 66886 72050 66938
rect 72102 66886 72114 66938
rect 72166 66886 74980 66938
rect 65320 66864 74980 66886
rect 63236 66484 63264 66792
rect 64874 66484 64880 66496
rect 63236 66456 64880 66484
rect 64874 66444 64880 66456
rect 64932 66444 64938 66496
rect 65320 66394 74980 66416
rect 65320 66342 74210 66394
rect 74262 66342 74274 66394
rect 74326 66342 74338 66394
rect 74390 66342 74402 66394
rect 74454 66342 74466 66394
rect 74518 66342 74980 66394
rect 65320 66320 74980 66342
rect 65320 65850 74980 65872
rect 63236 65668 63264 65816
rect 65320 65798 71858 65850
rect 71910 65798 71922 65850
rect 71974 65798 71986 65850
rect 72038 65798 72050 65850
rect 72102 65798 72114 65850
rect 72166 65798 74980 65850
rect 65320 65776 74980 65798
rect 65978 65668 65984 65680
rect 63236 65640 65984 65668
rect 65978 65628 65984 65640
rect 66036 65628 66042 65680
rect 63236 65396 63264 65564
rect 66070 65396 66076 65408
rect 63236 65368 66076 65396
rect 66070 65356 66076 65368
rect 66128 65356 66134 65408
rect 65320 65306 74980 65328
rect 65320 65254 74210 65306
rect 74262 65254 74274 65306
rect 74326 65254 74338 65306
rect 74390 65254 74402 65306
rect 74454 65254 74466 65306
rect 74518 65254 74980 65306
rect 65320 65232 74980 65254
rect 65320 64762 74980 64784
rect 65320 64710 71858 64762
rect 71910 64710 71922 64762
rect 71974 64710 71986 64762
rect 72038 64710 72050 64762
rect 72102 64710 72114 64762
rect 72166 64710 74980 64762
rect 65320 64688 74980 64710
rect 63236 64308 63264 64612
rect 64874 64308 64880 64320
rect 63236 64280 64880 64308
rect 64874 64268 64880 64280
rect 64932 64268 64938 64320
rect 65320 64218 74980 64240
rect 65320 64166 74210 64218
rect 74262 64166 74274 64218
rect 74326 64166 74338 64218
rect 74390 64166 74402 64218
rect 74454 64166 74466 64218
rect 74518 64166 74980 64218
rect 65320 64144 74980 64166
rect 65320 63674 74980 63696
rect 63236 63560 63264 63636
rect 65320 63622 71858 63674
rect 71910 63622 71922 63674
rect 71974 63622 71986 63674
rect 72038 63622 72050 63674
rect 72102 63622 72114 63674
rect 72166 63622 74980 63674
rect 65320 63600 74980 63622
rect 64966 63560 64972 63572
rect 63236 63532 64972 63560
rect 64966 63520 64972 63532
rect 65024 63520 65030 63572
rect 65702 63452 65708 63504
rect 65760 63452 65766 63504
rect 63236 63084 63264 63384
rect 66349 63359 66407 63365
rect 66349 63325 66361 63359
rect 66395 63356 66407 63359
rect 68002 63356 68008 63368
rect 66395 63328 68008 63356
rect 66395 63325 66407 63328
rect 66349 63319 66407 63325
rect 68002 63316 68008 63328
rect 68060 63316 68066 63368
rect 65320 63130 74980 63152
rect 63586 63084 63592 63096
rect 63236 63056 63592 63084
rect 63586 63044 63592 63056
rect 63644 63044 63650 63096
rect 65320 63078 74210 63130
rect 74262 63078 74274 63130
rect 74326 63078 74338 63130
rect 74390 63078 74402 63130
rect 74454 63078 74466 63130
rect 74518 63078 74980 63130
rect 65320 63056 74980 63078
rect 65320 62586 74980 62608
rect 65320 62534 71858 62586
rect 71910 62534 71922 62586
rect 71974 62534 71986 62586
rect 72038 62534 72050 62586
rect 72102 62534 72114 62586
rect 72166 62534 74980 62586
rect 65320 62512 74980 62534
rect 63236 62132 63264 62432
rect 64874 62132 64880 62144
rect 63236 62104 64880 62132
rect 64874 62092 64880 62104
rect 64932 62092 64938 62144
rect 65320 62042 74980 62064
rect 65320 61990 74210 62042
rect 74262 61990 74274 62042
rect 74326 61990 74338 62042
rect 74390 61990 74402 62042
rect 74454 61990 74466 62042
rect 74518 61990 74980 62042
rect 65320 61968 74980 61990
rect 65518 61888 65524 61940
rect 65576 61928 65582 61940
rect 65613 61931 65671 61937
rect 65613 61928 65625 61931
rect 65576 61900 65625 61928
rect 65576 61888 65582 61900
rect 65613 61897 65625 61900
rect 65659 61897 65671 61931
rect 65613 61891 65671 61897
rect 66257 61727 66315 61733
rect 66257 61693 66269 61727
rect 66303 61724 66315 61727
rect 66530 61724 66536 61736
rect 66303 61696 66536 61724
rect 66303 61693 66315 61696
rect 66257 61687 66315 61693
rect 66530 61684 66536 61696
rect 66588 61684 66594 61736
rect 65320 61498 74980 61520
rect 63236 61316 63264 61456
rect 65320 61446 71858 61498
rect 71910 61446 71922 61498
rect 71974 61446 71986 61498
rect 72038 61446 72050 61498
rect 72102 61446 72114 61498
rect 72166 61446 74980 61498
rect 65320 61424 74980 61446
rect 66162 61316 66168 61328
rect 63236 61288 66168 61316
rect 66162 61276 66168 61288
rect 66220 61276 66226 61328
rect 63494 61218 63500 61230
rect 63250 61190 63500 61218
rect 63494 61178 63500 61190
rect 63552 61178 63558 61230
rect 65320 60954 74980 60976
rect 65320 60902 74210 60954
rect 74262 60902 74274 60954
rect 74326 60902 74338 60954
rect 74390 60902 74402 60954
rect 74454 60902 74466 60954
rect 74518 60902 74980 60954
rect 65320 60880 74980 60902
rect 65320 60410 74980 60432
rect 65320 60358 71858 60410
rect 71910 60358 71922 60410
rect 71974 60358 71986 60410
rect 72038 60358 72050 60410
rect 72102 60358 72114 60410
rect 72166 60358 74980 60410
rect 65320 60336 74980 60358
rect 63144 60268 63816 60296
rect 63144 60252 63172 60268
rect 63788 60228 63816 60268
rect 65610 60256 65616 60308
rect 65668 60256 65674 60308
rect 64874 60228 64880 60240
rect 63788 60200 64880 60228
rect 64874 60188 64880 60200
rect 64932 60188 64938 60240
rect 66257 60095 66315 60101
rect 66257 60061 66269 60095
rect 66303 60092 66315 60095
rect 67082 60092 67088 60104
rect 66303 60064 67088 60092
rect 66303 60061 66315 60064
rect 66257 60055 66315 60061
rect 67082 60052 67088 60064
rect 67140 60052 67146 60104
rect 65320 59866 74980 59888
rect 65320 59814 74210 59866
rect 74262 59814 74274 59866
rect 74326 59814 74338 59866
rect 74390 59814 74402 59866
rect 74454 59814 74466 59866
rect 74518 59814 74980 59866
rect 65320 59792 74980 59814
rect 65320 59322 74980 59344
rect 63236 59140 63264 59276
rect 65320 59270 71858 59322
rect 71910 59270 71922 59322
rect 71974 59270 71986 59322
rect 72038 59270 72050 59322
rect 72102 59270 72114 59322
rect 72166 59270 74980 59322
rect 65320 59248 74980 59270
rect 65702 59140 65708 59152
rect 63236 59112 65708 59140
rect 65702 59100 65708 59112
rect 65760 59100 65766 59152
rect 71314 59072 71320 59084
rect 63236 59044 71320 59072
rect 63236 59024 63264 59044
rect 71314 59032 71320 59044
rect 71372 59032 71378 59084
rect 65320 58778 74980 58800
rect 65320 58726 74210 58778
rect 74262 58726 74274 58778
rect 74326 58726 74338 58778
rect 74390 58726 74402 58778
rect 74454 58726 74466 58778
rect 74518 58726 74980 58778
rect 65320 58704 74980 58726
rect 65334 58624 65340 58676
rect 65392 58664 65398 58676
rect 65613 58667 65671 58673
rect 65613 58664 65625 58667
rect 65392 58636 65625 58664
rect 65392 58624 65398 58636
rect 65613 58633 65625 58636
rect 65659 58633 65671 58667
rect 65613 58627 65671 58633
rect 66254 58420 66260 58472
rect 66312 58420 66318 58472
rect 65320 58234 74980 58256
rect 65320 58182 71858 58234
rect 71910 58182 71922 58234
rect 71974 58182 71986 58234
rect 72038 58182 72050 58234
rect 72102 58182 72114 58234
rect 72166 58182 74980 58234
rect 65320 58160 74980 58182
rect 63236 58052 63264 58072
rect 64874 58052 64880 58064
rect 63236 58024 64880 58052
rect 64874 58012 64880 58024
rect 64932 58012 64938 58064
rect 65320 57690 74980 57712
rect 65320 57638 74210 57690
rect 74262 57638 74274 57690
rect 74326 57638 74338 57690
rect 74390 57638 74402 57690
rect 74454 57638 74466 57690
rect 74518 57638 74980 57690
rect 65320 57616 74980 57638
rect 65320 57146 74980 57168
rect 63236 56964 63264 57096
rect 65320 57094 71858 57146
rect 71910 57094 71922 57146
rect 71974 57094 71986 57146
rect 72038 57094 72050 57146
rect 72102 57094 72114 57146
rect 72166 57094 74980 57146
rect 65320 57072 74980 57094
rect 65426 56992 65432 57044
rect 65484 57032 65490 57044
rect 65613 57035 65671 57041
rect 65613 57032 65625 57035
rect 65484 57004 65625 57032
rect 65484 56992 65490 57004
rect 65613 57001 65625 57004
rect 65659 57001 65671 57035
rect 65613 56995 65671 57001
rect 65518 56964 65524 56976
rect 63236 56936 65524 56964
rect 65518 56924 65524 56936
rect 65576 56924 65582 56976
rect 63236 56624 63264 56844
rect 66257 56831 66315 56837
rect 66257 56797 66269 56831
rect 66303 56828 66315 56831
rect 69290 56828 69296 56840
rect 66303 56800 69296 56828
rect 66303 56797 66315 56800
rect 66257 56791 66315 56797
rect 69290 56788 69296 56800
rect 69348 56788 69354 56840
rect 63678 56624 63684 56636
rect 63236 56596 63684 56624
rect 63678 56584 63684 56596
rect 63736 56584 63742 56636
rect 65320 56602 74980 56624
rect 65320 56550 74210 56602
rect 74262 56550 74274 56602
rect 74326 56550 74338 56602
rect 74390 56550 74402 56602
rect 74454 56550 74466 56602
rect 74518 56550 74980 56602
rect 65320 56528 74980 56550
rect 65320 56058 74980 56080
rect 65320 56006 71858 56058
rect 71910 56006 71922 56058
rect 71974 56006 71986 56058
rect 72038 56006 72050 56058
rect 72102 56006 72114 56058
rect 72166 56006 74980 56058
rect 65320 55984 74980 56006
rect 63236 55604 63264 55892
rect 64874 55604 64880 55616
rect 63236 55576 64880 55604
rect 64874 55564 64880 55576
rect 64932 55564 64938 55616
rect 65320 55514 74980 55536
rect 65320 55462 74210 55514
rect 74262 55462 74274 55514
rect 74326 55462 74338 55514
rect 74390 55462 74402 55514
rect 74454 55462 74466 55514
rect 74518 55462 74980 55514
rect 65320 55440 74980 55462
rect 65150 55360 65156 55412
rect 65208 55400 65214 55412
rect 65613 55403 65671 55409
rect 65613 55400 65625 55403
rect 65208 55372 65625 55400
rect 65208 55360 65214 55372
rect 65613 55369 65625 55372
rect 65659 55369 65671 55403
rect 65613 55363 65671 55369
rect 66257 55267 66315 55273
rect 66257 55233 66269 55267
rect 66303 55264 66315 55267
rect 69106 55264 69112 55276
rect 66303 55236 69112 55264
rect 66303 55233 66315 55236
rect 66257 55227 66315 55233
rect 69106 55224 69112 55236
rect 69164 55224 69170 55276
rect 65320 54970 74980 54992
rect 65320 54918 71858 54970
rect 71910 54918 71922 54970
rect 71974 54918 71986 54970
rect 72038 54918 72050 54970
rect 72102 54918 72114 54970
rect 72166 54918 74980 54970
rect 63236 54788 63264 54916
rect 65320 54896 74980 54918
rect 65334 54788 65340 54800
rect 63236 54760 65340 54788
rect 65334 54748 65340 54760
rect 65392 54748 65398 54800
rect 63144 54652 63172 54664
rect 71222 54652 71228 54664
rect 63144 54624 71228 54652
rect 71222 54612 71228 54624
rect 71280 54612 71286 54664
rect 65320 54426 74980 54448
rect 65320 54374 74210 54426
rect 74262 54374 74274 54426
rect 74326 54374 74338 54426
rect 74390 54374 74402 54426
rect 74454 54374 74466 54426
rect 74518 54374 74980 54426
rect 65320 54352 74980 54374
rect 65320 53882 74980 53904
rect 65320 53830 71858 53882
rect 71910 53830 71922 53882
rect 71974 53830 71986 53882
rect 72038 53830 72050 53882
rect 72102 53830 72114 53882
rect 72166 53830 74980 53882
rect 65320 53808 74980 53830
rect 63236 53564 63264 53712
rect 65794 53592 65800 53644
rect 65852 53592 65858 53644
rect 64874 53564 64880 53576
rect 63236 53536 64880 53564
rect 64874 53524 64880 53536
rect 64932 53524 64938 53576
rect 66993 53567 67051 53573
rect 66993 53533 67005 53567
rect 67039 53564 67051 53567
rect 69382 53564 69388 53576
rect 67039 53536 69388 53564
rect 67039 53533 67051 53536
rect 66993 53527 67051 53533
rect 69382 53524 69388 53536
rect 69440 53524 69446 53576
rect 63236 53428 63264 53432
rect 69014 53428 69020 53440
rect 63236 53400 69020 53428
rect 69014 53388 69020 53400
rect 69072 53388 69078 53440
rect 65320 53338 74980 53360
rect 65320 53286 74210 53338
rect 74262 53286 74274 53338
rect 74326 53286 74338 53338
rect 74390 53286 74402 53338
rect 74454 53286 74466 53338
rect 74518 53286 74980 53338
rect 65320 53264 74980 53286
rect 65242 53184 65248 53236
rect 65300 53224 65306 53236
rect 65613 53227 65671 53233
rect 65613 53224 65625 53227
rect 65300 53196 65625 53224
rect 65300 53184 65306 53196
rect 65613 53193 65625 53196
rect 65659 53193 65671 53227
rect 65613 53187 65671 53193
rect 66257 53023 66315 53029
rect 66257 52989 66269 53023
rect 66303 53020 66315 53023
rect 66346 53020 66352 53032
rect 66303 52992 66352 53020
rect 66303 52989 66315 52992
rect 66257 52983 66315 52989
rect 66346 52980 66352 52992
rect 66404 52980 66410 53032
rect 65320 52794 74980 52816
rect 65320 52742 71858 52794
rect 71910 52742 71922 52794
rect 71974 52742 71986 52794
rect 72038 52742 72050 52794
rect 72102 52742 72114 52794
rect 72166 52742 74980 52794
rect 63236 52612 63264 52736
rect 65320 52720 74980 52742
rect 65426 52612 65432 52624
rect 63236 52584 65432 52612
rect 65426 52572 65432 52584
rect 65484 52572 65490 52624
rect 63236 52476 63264 52484
rect 63770 52476 63776 52488
rect 63236 52448 63776 52476
rect 63770 52436 63776 52448
rect 63828 52436 63834 52488
rect 65610 52436 65616 52488
rect 65668 52436 65674 52488
rect 65889 52479 65947 52485
rect 65889 52445 65901 52479
rect 65935 52445 65947 52479
rect 65889 52439 65947 52445
rect 65904 52408 65932 52439
rect 63236 52380 65932 52408
rect 63236 52171 63264 52380
rect 65320 52250 74980 52272
rect 65320 52198 74210 52250
rect 74262 52198 74274 52250
rect 74326 52198 74338 52250
rect 74390 52198 74402 52250
rect 74454 52198 74466 52250
rect 74518 52198 74980 52250
rect 65320 52176 74980 52198
rect 65610 52136 65616 52148
rect 63604 52108 65616 52136
rect 63250 52080 63632 52108
rect 65610 52096 65616 52108
rect 65668 52096 65674 52148
rect 65058 51960 65064 52012
rect 65116 52000 65122 52012
rect 65613 52003 65671 52009
rect 65613 52000 65625 52003
rect 65116 51972 65625 52000
rect 65116 51960 65122 51972
rect 65613 51969 65625 51972
rect 65659 51969 65671 52003
rect 65613 51963 65671 51969
rect 66257 51935 66315 51941
rect 66257 51901 66269 51935
rect 66303 51932 66315 51935
rect 67542 51932 67548 51944
rect 66303 51904 67548 51932
rect 66303 51901 66315 51904
rect 66257 51895 66315 51901
rect 67542 51892 67548 51904
rect 67600 51892 67606 51944
rect 65320 51706 74980 51728
rect 65320 51654 71858 51706
rect 71910 51654 71922 51706
rect 71974 51654 71986 51706
rect 72038 51654 72050 51706
rect 72102 51654 72114 51706
rect 72166 51654 74980 51706
rect 65320 51632 74980 51654
rect 63236 51524 63264 51532
rect 64874 51524 64880 51536
rect 63236 51496 64880 51524
rect 64874 51484 64880 51496
rect 64932 51524 64938 51536
rect 65794 51524 65800 51536
rect 64932 51496 65800 51524
rect 64932 51484 64938 51496
rect 65794 51484 65800 51496
rect 65852 51484 65858 51536
rect 65320 51162 74980 51184
rect 65320 51110 74210 51162
rect 74262 51110 74274 51162
rect 74326 51110 74338 51162
rect 74390 51110 74402 51162
rect 74454 51110 74466 51162
rect 74518 51110 74980 51162
rect 65320 51088 74980 51110
rect 65320 50618 74980 50640
rect 65320 50566 71858 50618
rect 71910 50566 71922 50618
rect 71974 50566 71986 50618
rect 72038 50566 72050 50618
rect 72102 50566 72114 50618
rect 72166 50566 74980 50618
rect 63236 50436 63264 50556
rect 65320 50544 74980 50566
rect 65613 50507 65671 50513
rect 65613 50473 65625 50507
rect 65659 50504 65671 50507
rect 65978 50504 65984 50516
rect 65659 50476 65984 50504
rect 65659 50473 65671 50476
rect 65613 50467 65671 50473
rect 65978 50464 65984 50476
rect 66036 50464 66042 50516
rect 65150 50436 65156 50448
rect 63236 50408 65156 50436
rect 65150 50396 65156 50408
rect 65208 50396 65214 50448
rect 66257 50371 66315 50377
rect 66257 50337 66269 50371
rect 66303 50368 66315 50371
rect 67634 50368 67640 50380
rect 66303 50340 67640 50368
rect 66303 50337 66315 50340
rect 66257 50331 66315 50337
rect 67634 50328 67640 50340
rect 67692 50328 67698 50380
rect 63236 50300 63264 50304
rect 63862 50300 63868 50312
rect 63236 50272 63868 50300
rect 63862 50260 63868 50272
rect 63920 50260 63926 50312
rect 66349 50303 66407 50309
rect 66349 50269 66361 50303
rect 66395 50269 66407 50303
rect 66349 50263 66407 50269
rect 66364 50232 66392 50263
rect 63236 50204 66392 50232
rect 63236 49996 63264 50204
rect 65320 50074 74980 50096
rect 65320 50022 74210 50074
rect 74262 50022 74274 50074
rect 74326 50022 74338 50074
rect 74390 50022 74402 50074
rect 74454 50022 74466 50074
rect 74518 50022 74980 50074
rect 65320 50000 74980 50022
rect 63144 49552 63172 49657
rect 65613 49623 65671 49629
rect 65613 49620 65625 49623
rect 63420 49592 65625 49620
rect 63420 49552 63448 49592
rect 65613 49589 65625 49592
rect 65659 49589 65671 49623
rect 65613 49583 65671 49589
rect 63144 49524 63448 49552
rect 65320 49530 74980 49552
rect 65320 49478 71858 49530
rect 71910 49478 71922 49530
rect 71974 49478 71986 49530
rect 72038 49478 72050 49530
rect 72102 49478 72114 49530
rect 72166 49478 74980 49530
rect 65320 49456 74980 49478
rect 63402 49172 63408 49224
rect 63460 49212 63466 49224
rect 65613 49215 65671 49221
rect 65613 49212 65625 49215
rect 63460 49184 65625 49212
rect 63460 49172 63466 49184
rect 65613 49181 65625 49184
rect 65659 49181 65671 49215
rect 65613 49175 65671 49181
rect 65320 48986 74980 49008
rect 65320 48934 74210 48986
rect 74262 48934 74274 48986
rect 74326 48934 74338 48986
rect 74390 48934 74402 48986
rect 74454 48934 74466 48986
rect 74518 48934 74980 48986
rect 65320 48912 74980 48934
rect 64966 48832 64972 48884
rect 65024 48872 65030 48884
rect 65613 48875 65671 48881
rect 65613 48872 65625 48875
rect 65024 48844 65625 48872
rect 65024 48832 65030 48844
rect 65613 48841 65625 48844
rect 65659 48841 65671 48875
rect 65613 48835 65671 48841
rect 63250 48804 63540 48809
rect 69750 48804 69756 48816
rect 63250 48781 69756 48804
rect 63512 48776 69756 48781
rect 69750 48764 69756 48776
rect 69808 48764 69814 48816
rect 63402 48729 63408 48741
rect 63250 48701 63408 48729
rect 63402 48689 63408 48701
rect 63460 48689 63466 48741
rect 66257 48671 66315 48677
rect 66257 48637 66269 48671
rect 66303 48668 66315 48671
rect 69566 48668 69572 48680
rect 66303 48640 69572 48668
rect 66303 48637 66315 48640
rect 66257 48631 66315 48637
rect 69566 48628 69572 48640
rect 69624 48628 69630 48680
rect 65320 48442 74980 48464
rect 65320 48390 71858 48442
rect 71910 48390 71922 48442
rect 71974 48390 71986 48442
rect 72038 48390 72050 48442
rect 72102 48390 72114 48442
rect 72166 48390 74980 48442
rect 65320 48368 74980 48390
rect 69198 48124 69204 48136
rect 63236 48096 69204 48124
rect 63236 48087 63264 48096
rect 69198 48084 69204 48096
rect 69256 48084 69262 48136
rect 63236 47716 63264 48007
rect 65320 47898 74980 47920
rect 65320 47846 74210 47898
rect 74262 47846 74274 47898
rect 74326 47846 74338 47898
rect 74390 47846 74402 47898
rect 74454 47846 74466 47898
rect 74518 47846 74980 47898
rect 65320 47824 74980 47846
rect 64966 47716 64972 47728
rect 63236 47688 64972 47716
rect 64966 47676 64972 47688
rect 65024 47676 65030 47728
rect 63250 47376 63632 47393
rect 64874 47376 64880 47388
rect 63250 47365 64880 47376
rect 63604 47348 64880 47365
rect 64874 47336 64880 47348
rect 64932 47336 64938 47388
rect 65320 47354 74980 47376
rect 63402 47313 63408 47325
rect 63250 47285 63408 47313
rect 63402 47273 63408 47285
rect 63460 47273 63466 47325
rect 65320 47302 71858 47354
rect 71910 47302 71922 47354
rect 71974 47302 71986 47354
rect 72038 47302 72050 47354
rect 72102 47302 72114 47354
rect 72166 47302 74980 47354
rect 65320 47280 74980 47302
rect 65613 47243 65671 47249
rect 65613 47209 65625 47243
rect 65659 47240 65671 47243
rect 66162 47240 66168 47252
rect 65659 47212 66168 47240
rect 65659 47209 65671 47212
rect 65613 47203 65671 47209
rect 66162 47200 66168 47212
rect 66220 47200 66226 47252
rect 66349 47107 66407 47113
rect 66349 47073 66361 47107
rect 66395 47104 66407 47107
rect 70762 47104 70768 47116
rect 66395 47076 70768 47104
rect 66395 47073 66407 47076
rect 66349 47067 66407 47073
rect 70762 47064 70768 47076
rect 70820 47064 70826 47116
rect 66257 47039 66315 47045
rect 66257 47005 66269 47039
rect 66303 47036 66315 47039
rect 69658 47036 69664 47048
rect 66303 47008 69664 47036
rect 66303 47005 66315 47008
rect 66257 46999 66315 47005
rect 69658 46996 69664 47008
rect 69716 46996 69722 47048
rect 66622 46928 66628 46980
rect 66680 46928 66686 46980
rect 65320 46810 74980 46832
rect 65320 46758 74210 46810
rect 74262 46758 74274 46810
rect 74326 46758 74338 46810
rect 74390 46758 74402 46810
rect 74454 46758 74466 46810
rect 74518 46758 74980 46810
rect 65320 46736 74980 46758
rect 65320 46266 74980 46288
rect 65320 46214 71858 46266
rect 71910 46214 71922 46266
rect 71974 46214 71986 46266
rect 72038 46214 72050 46266
rect 72102 46214 72114 46266
rect 72166 46214 74980 46266
rect 65320 46192 74980 46214
rect 63250 45949 63632 45977
rect 63604 45948 63632 45949
rect 65058 45948 65064 45960
rect 63604 45920 65064 45948
rect 65058 45908 65064 45920
rect 65116 45908 65122 45960
rect 63236 45608 63264 45883
rect 65320 45722 74980 45744
rect 65320 45670 74210 45722
rect 74262 45670 74274 45722
rect 74326 45670 74338 45722
rect 74390 45670 74402 45722
rect 74454 45670 74466 45722
rect 74518 45670 74980 45722
rect 65320 45648 74980 45670
rect 66990 45608 66996 45620
rect 63236 45580 66996 45608
rect 66990 45568 66996 45580
rect 67048 45568 67054 45620
rect 65610 45500 65616 45552
rect 65668 45500 65674 45552
rect 66257 45407 66315 45413
rect 66257 45373 66269 45407
rect 66303 45404 66315 45407
rect 67174 45404 67180 45416
rect 66303 45376 67180 45404
rect 66303 45373 66315 45376
rect 66257 45367 66315 45373
rect 67174 45364 67180 45376
rect 67232 45364 67238 45416
rect 63250 45268 63632 45269
rect 67266 45268 67272 45280
rect 63250 45241 67272 45268
rect 63604 45240 67272 45241
rect 67266 45228 67272 45240
rect 67324 45228 67330 45280
rect 65320 45178 74980 45200
rect 63236 44860 63264 45175
rect 65320 45126 71858 45178
rect 71910 45126 71922 45178
rect 71974 45126 71986 45178
rect 72038 45126 72050 45178
rect 72102 45126 72114 45178
rect 72166 45126 74980 45178
rect 65320 45104 74980 45126
rect 66806 44860 66812 44872
rect 63236 44832 66812 44860
rect 66806 44820 66812 44832
rect 66864 44820 66870 44872
rect 64966 44684 64972 44736
rect 65024 44724 65030 44736
rect 65610 44724 65616 44736
rect 65024 44696 65616 44724
rect 65024 44684 65030 44696
rect 65610 44684 65616 44696
rect 65668 44684 65674 44736
rect 65320 44634 74980 44656
rect 64966 44588 64972 44600
rect 63236 44560 64972 44588
rect 63236 44547 63264 44560
rect 64966 44548 64972 44560
rect 65024 44548 65030 44600
rect 65320 44582 74210 44634
rect 74262 44582 74274 44634
rect 74326 44582 74338 44634
rect 74390 44582 74402 44634
rect 74454 44582 74466 44634
rect 74518 44582 74980 44634
rect 65320 44560 74980 44582
rect 63236 44180 63264 44467
rect 65794 44180 65800 44192
rect 63236 44152 65800 44180
rect 65794 44140 65800 44152
rect 65852 44140 65858 44192
rect 66622 44140 66628 44192
rect 66680 44180 66686 44192
rect 70854 44180 70860 44192
rect 66680 44152 70860 44180
rect 66680 44140 66686 44152
rect 70854 44140 70860 44152
rect 70912 44140 70918 44192
rect 65320 44090 74980 44112
rect 65320 44038 71858 44090
rect 71910 44038 71922 44090
rect 71974 44038 71986 44090
rect 72038 44038 72050 44090
rect 72102 44038 72114 44090
rect 72166 44038 74980 44090
rect 65320 44016 74980 44038
rect 65518 43936 65524 43988
rect 65576 43976 65582 43988
rect 65613 43979 65671 43985
rect 65613 43976 65625 43979
rect 65576 43948 65625 43976
rect 65576 43936 65582 43948
rect 65613 43945 65625 43948
rect 65659 43945 65671 43979
rect 65613 43939 65671 43945
rect 66257 43843 66315 43849
rect 63236 43772 63264 43839
rect 66257 43809 66269 43843
rect 66303 43840 66315 43843
rect 66438 43840 66444 43852
rect 66303 43812 66444 43840
rect 66303 43809 66315 43812
rect 66257 43803 66315 43809
rect 66438 43800 66444 43812
rect 66496 43800 66502 43852
rect 65978 43772 65984 43784
rect 63236 43744 65984 43772
rect 65978 43732 65984 43744
rect 66036 43732 66042 43784
rect 66349 43775 66407 43781
rect 66349 43741 66361 43775
rect 66395 43741 66407 43775
rect 66349 43735 66407 43741
rect 66364 43704 66392 43735
rect 63236 43676 66392 43704
rect 63236 43654 63264 43676
rect 65320 43546 74980 43568
rect 65320 43494 74210 43546
rect 74262 43494 74274 43546
rect 74326 43494 74338 43546
rect 74390 43494 74402 43546
rect 74454 43494 74466 43546
rect 74518 43494 74980 43546
rect 65320 43472 74980 43494
rect 63236 43160 63264 43270
rect 63954 43160 63960 43172
rect 63236 43132 63960 43160
rect 63954 43120 63960 43132
rect 64012 43120 64018 43172
rect 63236 42820 63264 43018
rect 65320 43002 74980 43024
rect 65320 42950 71858 43002
rect 71910 42950 71922 43002
rect 71974 42950 71986 43002
rect 72038 42950 72050 43002
rect 72102 42950 72114 43002
rect 72166 42950 74980 43002
rect 65320 42928 74980 42950
rect 66162 42820 66168 42832
rect 63236 42792 66168 42820
rect 66162 42780 66168 42792
rect 66220 42780 66226 42832
rect 68002 42712 68008 42764
rect 68060 42712 68066 42764
rect 65613 42687 65671 42693
rect 65613 42684 65625 42687
rect 63236 42656 65625 42684
rect 63236 42402 63264 42656
rect 65613 42653 65625 42656
rect 65659 42653 65671 42687
rect 65613 42647 65671 42653
rect 68649 42687 68707 42693
rect 68649 42653 68661 42687
rect 68695 42684 68707 42687
rect 70118 42684 70124 42696
rect 68695 42656 70124 42684
rect 68695 42653 68707 42656
rect 68649 42647 68707 42653
rect 70118 42644 70124 42656
rect 70176 42644 70182 42696
rect 65320 42458 74980 42480
rect 65320 42406 74210 42458
rect 74262 42406 74274 42458
rect 74326 42406 74338 42458
rect 74390 42406 74402 42458
rect 74454 42406 74466 42458
rect 74518 42406 74980 42458
rect 65320 42384 74980 42406
rect 65334 42304 65340 42356
rect 65392 42344 65398 42356
rect 65613 42347 65671 42353
rect 65613 42344 65625 42347
rect 65392 42316 65625 42344
rect 65392 42304 65398 42316
rect 65613 42313 65625 42316
rect 65659 42313 65671 42347
rect 65613 42307 65671 42313
rect 66257 42143 66315 42149
rect 66257 42109 66269 42143
rect 66303 42140 66315 42143
rect 66714 42140 66720 42152
rect 66303 42112 66720 42140
rect 66303 42109 66315 42112
rect 66257 42103 66315 42109
rect 66714 42100 66720 42112
rect 66772 42100 66778 42152
rect 65426 42072 65432 42084
rect 65260 42044 65432 42072
rect 63236 41732 63264 42042
rect 65260 41800 65288 42044
rect 65426 42032 65432 42044
rect 65484 42032 65490 42084
rect 65320 41914 74980 41936
rect 65320 41862 71858 41914
rect 71910 41862 71922 41914
rect 71974 41862 71986 41914
rect 72038 41862 72050 41914
rect 72102 41862 72114 41914
rect 72166 41862 74980 41914
rect 65320 41840 74980 41862
rect 65426 41800 65432 41812
rect 65260 41772 65432 41800
rect 65426 41760 65432 41772
rect 65484 41760 65490 41812
rect 66530 41760 66536 41812
rect 66588 41800 66594 41812
rect 66717 41803 66775 41809
rect 66717 41800 66729 41803
rect 66588 41772 66729 41800
rect 66588 41760 66594 41772
rect 66717 41769 66729 41772
rect 66763 41769 66775 41803
rect 66717 41763 66775 41769
rect 65150 41732 65156 41744
rect 63236 41704 65156 41732
rect 65150 41692 65156 41704
rect 65208 41692 65214 41744
rect 67361 41599 67419 41605
rect 67361 41565 67373 41599
rect 67407 41596 67419 41599
rect 68554 41596 68560 41608
rect 67407 41568 68560 41596
rect 67407 41565 67419 41568
rect 67361 41559 67419 41565
rect 68554 41556 68560 41568
rect 68612 41556 68618 41608
rect 65320 41370 74980 41392
rect 65320 41318 74210 41370
rect 74262 41318 74274 41370
rect 74326 41318 74338 41370
rect 74390 41318 74402 41370
rect 74454 41318 74466 41370
rect 74518 41318 74980 41370
rect 65320 41296 74980 41318
rect 63236 40984 63264 41090
rect 64046 40984 64052 40996
rect 63236 40956 64052 40984
rect 64046 40944 64052 40956
rect 64104 40944 64110 40996
rect 65794 40876 65800 40928
rect 65852 40876 65858 40928
rect 63236 40576 63264 40838
rect 65320 40826 74980 40848
rect 65320 40774 71858 40826
rect 71910 40774 71922 40826
rect 71974 40774 71986 40826
rect 72038 40774 72050 40826
rect 72102 40774 72114 40826
rect 72166 40774 74980 40826
rect 65320 40752 74980 40774
rect 67082 40672 67088 40724
rect 67140 40672 67146 40724
rect 65334 40576 65340 40588
rect 63236 40548 65340 40576
rect 65334 40536 65340 40548
rect 65392 40536 65398 40588
rect 65702 40536 65708 40588
rect 65760 40576 65766 40588
rect 65797 40579 65855 40585
rect 65797 40576 65809 40579
rect 65760 40548 65809 40576
rect 65760 40536 65766 40548
rect 65797 40545 65809 40548
rect 65843 40545 65855 40579
rect 65797 40539 65855 40545
rect 66530 40468 66536 40520
rect 66588 40508 66594 40520
rect 66809 40511 66867 40517
rect 66809 40508 66821 40511
rect 66588 40480 66821 40508
rect 66588 40468 66594 40480
rect 66809 40477 66821 40480
rect 66855 40477 66867 40511
rect 66809 40471 66867 40477
rect 67729 40511 67787 40517
rect 67729 40477 67741 40511
rect 67775 40508 67787 40511
rect 68186 40508 68192 40520
rect 67775 40480 68192 40508
rect 67775 40477 67787 40480
rect 67729 40471 67787 40477
rect 68186 40468 68192 40480
rect 68244 40468 68250 40520
rect 65702 40332 65708 40384
rect 65760 40372 65766 40384
rect 65978 40372 65984 40384
rect 65760 40344 65984 40372
rect 65760 40332 65766 40344
rect 65978 40332 65984 40344
rect 66036 40332 66042 40384
rect 65320 40282 74980 40304
rect 65320 40230 74210 40282
rect 74262 40230 74274 40282
rect 74326 40230 74338 40282
rect 74390 40230 74402 40282
rect 74454 40230 74466 40282
rect 74518 40230 74980 40282
rect 65320 40208 74980 40230
rect 65426 40128 65432 40180
rect 65484 40168 65490 40180
rect 65613 40171 65671 40177
rect 65613 40168 65625 40171
rect 65484 40140 65625 40168
rect 65484 40128 65490 40140
rect 65613 40137 65625 40140
rect 65659 40137 65671 40171
rect 65613 40131 65671 40137
rect 66257 39967 66315 39973
rect 66257 39933 66269 39967
rect 66303 39964 66315 39967
rect 66622 39964 66628 39976
rect 66303 39936 66628 39964
rect 66303 39933 66315 39936
rect 66257 39927 66315 39933
rect 66622 39924 66628 39936
rect 66680 39924 66686 39976
rect 63144 39868 63816 39896
rect 63144 39862 63172 39868
rect 63788 39828 63816 39868
rect 65150 39828 65156 39840
rect 63788 39800 65156 39828
rect 65150 39788 65156 39800
rect 65208 39788 65214 39840
rect 65320 39738 74980 39760
rect 65320 39686 71858 39738
rect 71910 39686 71922 39738
rect 71974 39686 71986 39738
rect 72038 39686 72050 39738
rect 72102 39686 72114 39738
rect 72166 39686 74980 39738
rect 65320 39664 74980 39686
rect 63402 39584 63408 39636
rect 63460 39624 63466 39636
rect 65518 39624 65524 39636
rect 63460 39596 65524 39624
rect 63460 39584 63466 39596
rect 65518 39584 65524 39596
rect 65576 39584 65582 39636
rect 65613 39627 65671 39633
rect 65613 39593 65625 39627
rect 65659 39624 65671 39627
rect 66254 39624 66260 39636
rect 65659 39596 66260 39624
rect 65659 39593 65671 39596
rect 65613 39587 65671 39593
rect 66254 39584 66260 39596
rect 66312 39584 66318 39636
rect 66257 39423 66315 39429
rect 66257 39389 66269 39423
rect 66303 39420 66315 39423
rect 67542 39420 67548 39432
rect 66303 39392 67548 39420
rect 66303 39389 66315 39392
rect 66257 39383 66315 39389
rect 67542 39380 67548 39392
rect 67600 39380 67606 39432
rect 65320 39194 74980 39216
rect 65320 39142 74210 39194
rect 74262 39142 74274 39194
rect 74326 39142 74338 39194
rect 74390 39142 74402 39194
rect 74454 39142 74466 39194
rect 74518 39142 74980 39194
rect 65320 39120 74980 39142
rect 65242 39040 65248 39092
rect 65300 39080 65306 39092
rect 65613 39083 65671 39089
rect 65613 39080 65625 39083
rect 65300 39052 65625 39080
rect 65300 39040 65306 39052
rect 65613 39049 65625 39052
rect 65659 39049 65671 39083
rect 65613 39043 65671 39049
rect 63402 38924 63408 38936
rect 63250 38896 63408 38924
rect 63402 38884 63408 38896
rect 63460 38884 63466 38936
rect 66257 38879 66315 38885
rect 66257 38845 66269 38879
rect 66303 38876 66315 38879
rect 69842 38876 69848 38888
rect 66303 38848 69848 38876
rect 66303 38845 66315 38848
rect 66257 38839 66315 38845
rect 69842 38836 69848 38848
rect 69900 38836 69906 38888
rect 65426 38740 65432 38752
rect 63236 38712 65432 38740
rect 63236 38658 63264 38712
rect 65426 38700 65432 38712
rect 65484 38700 65490 38752
rect 65320 38650 74980 38672
rect 65320 38598 71858 38650
rect 71910 38598 71922 38650
rect 71974 38598 71986 38650
rect 72038 38598 72050 38650
rect 72102 38598 72114 38650
rect 72166 38598 74980 38650
rect 65320 38576 74980 38598
rect 65613 38539 65671 38545
rect 65613 38505 65625 38539
rect 65659 38536 65671 38539
rect 69290 38536 69296 38548
rect 65659 38508 69296 38536
rect 65659 38505 65671 38508
rect 65613 38499 65671 38505
rect 69290 38496 69296 38508
rect 69348 38496 69354 38548
rect 65978 38428 65984 38480
rect 66036 38468 66042 38480
rect 66254 38468 66260 38480
rect 66036 38440 66260 38468
rect 66036 38428 66042 38440
rect 66254 38428 66260 38440
rect 66312 38428 66318 38480
rect 66257 38335 66315 38341
rect 66257 38301 66269 38335
rect 66303 38332 66315 38335
rect 69474 38332 69480 38344
rect 66303 38304 69480 38332
rect 66303 38301 66315 38304
rect 66257 38295 66315 38301
rect 69474 38292 69480 38304
rect 69532 38292 69538 38344
rect 65320 38106 74980 38128
rect 65320 38054 74210 38106
rect 74262 38054 74274 38106
rect 74326 38054 74338 38106
rect 74390 38054 74402 38106
rect 74454 38054 74466 38106
rect 74518 38054 74980 38106
rect 65320 38032 74980 38054
rect 66257 37995 66315 38001
rect 66257 37961 66269 37995
rect 66303 37992 66315 37995
rect 69106 37992 69112 38004
rect 66303 37964 69112 37992
rect 66303 37961 66315 37964
rect 66257 37955 66315 37961
rect 69106 37952 69112 37964
rect 69164 37952 69170 38004
rect 65705 37791 65763 37797
rect 65705 37757 65717 37791
rect 65751 37788 65763 37791
rect 70026 37788 70032 37800
rect 65751 37760 70032 37788
rect 65751 37757 65763 37760
rect 65705 37751 65763 37757
rect 70026 37748 70032 37760
rect 70084 37748 70090 37800
rect 63236 37380 63264 37682
rect 65320 37562 74980 37584
rect 65320 37510 71858 37562
rect 71910 37510 71922 37562
rect 71974 37510 71986 37562
rect 72038 37510 72050 37562
rect 72102 37510 72114 37562
rect 72166 37510 74980 37562
rect 65320 37488 74980 37510
rect 65150 37380 65156 37392
rect 63236 37352 65156 37380
rect 65150 37340 65156 37352
rect 65208 37340 65214 37392
rect 65610 37204 65616 37256
rect 65668 37204 65674 37256
rect 66257 37247 66315 37253
rect 66257 37213 66269 37247
rect 66303 37244 66315 37247
rect 67450 37244 67456 37256
rect 66303 37216 67456 37244
rect 66303 37213 66315 37216
rect 66257 37207 66315 37213
rect 67450 37204 67456 37216
rect 67508 37204 67514 37256
rect 65320 37018 74980 37040
rect 65320 36966 74210 37018
rect 74262 36966 74274 37018
rect 74326 36966 74338 37018
rect 74390 36966 74402 37018
rect 74454 36966 74466 37018
rect 74518 36966 74980 37018
rect 65320 36944 74980 36966
rect 65518 36864 65524 36916
rect 65576 36904 65582 36916
rect 65613 36907 65671 36913
rect 65613 36904 65625 36907
rect 65576 36876 65625 36904
rect 65576 36864 65582 36876
rect 65613 36873 65625 36876
rect 65659 36873 65671 36907
rect 65613 36867 65671 36873
rect 63236 36564 63264 36730
rect 64966 36728 64972 36780
rect 65024 36768 65030 36780
rect 65518 36768 65524 36780
rect 65024 36740 65524 36768
rect 65024 36728 65030 36740
rect 65518 36728 65524 36740
rect 65576 36728 65582 36780
rect 66257 36703 66315 36709
rect 66257 36669 66269 36703
rect 66303 36700 66315 36703
rect 66898 36700 66904 36712
rect 66303 36672 66904 36700
rect 66303 36669 66315 36672
rect 66257 36663 66315 36669
rect 66898 36660 66904 36672
rect 66956 36660 66962 36712
rect 64966 36564 64972 36576
rect 63236 36536 64972 36564
rect 64966 36524 64972 36536
rect 65024 36524 65030 36576
rect 63236 36156 63264 36478
rect 65320 36474 74980 36496
rect 65320 36422 71858 36474
rect 71910 36422 71922 36474
rect 71974 36422 71986 36474
rect 72038 36422 72050 36474
rect 72102 36422 72114 36474
rect 72166 36422 74980 36474
rect 65320 36400 74980 36422
rect 64874 36320 64880 36372
rect 64932 36360 64938 36372
rect 65613 36363 65671 36369
rect 65613 36360 65625 36363
rect 64932 36332 65625 36360
rect 64932 36320 64938 36332
rect 65613 36329 65625 36332
rect 65659 36329 65671 36363
rect 65613 36323 65671 36329
rect 66346 36320 66352 36372
rect 66404 36320 66410 36372
rect 66257 36227 66315 36233
rect 66257 36193 66269 36227
rect 66303 36224 66315 36227
rect 67358 36224 67364 36236
rect 66303 36196 67364 36224
rect 66303 36193 66315 36196
rect 66257 36187 66315 36193
rect 67358 36184 67364 36196
rect 67416 36184 67422 36236
rect 65978 36156 65984 36168
rect 63236 36128 65984 36156
rect 65978 36116 65984 36128
rect 66036 36116 66042 36168
rect 66993 36159 67051 36165
rect 66993 36125 67005 36159
rect 67039 36156 67051 36159
rect 68278 36156 68284 36168
rect 67039 36128 68284 36156
rect 67039 36125 67051 36128
rect 66993 36119 67051 36125
rect 68278 36116 68284 36128
rect 68336 36116 68342 36168
rect 65320 35930 74980 35952
rect 65320 35878 74210 35930
rect 74262 35878 74274 35930
rect 74326 35878 74338 35930
rect 74390 35878 74402 35930
rect 74454 35878 74466 35930
rect 74518 35878 74980 35930
rect 65320 35856 74980 35878
rect 66990 35776 66996 35828
rect 67048 35816 67054 35828
rect 67085 35819 67143 35825
rect 67085 35816 67097 35819
rect 67048 35788 67097 35816
rect 67048 35776 67054 35788
rect 67085 35785 67097 35788
rect 67131 35785 67143 35819
rect 67085 35779 67143 35785
rect 66809 35751 66867 35757
rect 66809 35717 66821 35751
rect 66855 35748 66867 35751
rect 69382 35748 69388 35760
rect 66855 35720 69388 35748
rect 66855 35717 66867 35720
rect 66809 35711 66867 35717
rect 69382 35708 69388 35720
rect 69440 35708 69446 35760
rect 64138 35640 64144 35692
rect 64196 35680 64202 35692
rect 65613 35683 65671 35689
rect 65613 35680 65625 35683
rect 64196 35652 65625 35680
rect 64196 35640 64202 35652
rect 65613 35649 65625 35652
rect 65659 35649 65671 35683
rect 65613 35643 65671 35649
rect 67729 35615 67787 35621
rect 67729 35581 67741 35615
rect 67775 35612 67787 35615
rect 68370 35612 68376 35624
rect 67775 35584 68376 35612
rect 67775 35581 67787 35584
rect 67729 35575 67787 35581
rect 68370 35572 68376 35584
rect 68428 35572 68434 35624
rect 63236 35204 63264 35502
rect 65320 35386 74980 35408
rect 65320 35334 71858 35386
rect 71910 35334 71922 35386
rect 71974 35334 71986 35386
rect 72038 35334 72050 35386
rect 72102 35334 72114 35386
rect 72166 35334 74980 35386
rect 65320 35312 74980 35334
rect 67910 35232 67916 35284
rect 67968 35272 67974 35284
rect 68005 35275 68063 35281
rect 68005 35272 68017 35275
rect 67968 35244 68017 35272
rect 67968 35232 67974 35244
rect 68005 35241 68017 35244
rect 68051 35241 68063 35275
rect 68005 35235 68063 35241
rect 64874 35204 64880 35216
rect 63236 35176 64880 35204
rect 64874 35164 64880 35176
rect 64932 35204 64938 35216
rect 65150 35204 65156 35216
rect 64932 35176 65156 35204
rect 64932 35164 64938 35176
rect 65150 35164 65156 35176
rect 65208 35164 65214 35216
rect 67361 35139 67419 35145
rect 67361 35105 67373 35139
rect 67407 35136 67419 35139
rect 69014 35136 69020 35148
rect 67407 35108 69020 35136
rect 67407 35105 67419 35108
rect 67361 35099 67419 35105
rect 69014 35096 69020 35108
rect 69072 35096 69078 35148
rect 68462 35028 68468 35080
rect 68520 35068 68526 35080
rect 68557 35071 68615 35077
rect 68557 35068 68569 35071
rect 68520 35040 68569 35068
rect 68520 35028 68526 35040
rect 68557 35037 68569 35040
rect 68603 35037 68615 35071
rect 68557 35031 68615 35037
rect 65610 34960 65616 35012
rect 65668 34960 65674 35012
rect 65320 34842 74980 34864
rect 65320 34790 74210 34842
rect 74262 34790 74274 34842
rect 74326 34790 74338 34842
rect 74390 34790 74402 34842
rect 74454 34790 74466 34842
rect 74518 34790 74980 34842
rect 65320 34768 74980 34790
rect 65058 34688 65064 34740
rect 65116 34728 65122 34740
rect 65613 34731 65671 34737
rect 65613 34728 65625 34731
rect 65116 34700 65625 34728
rect 65116 34688 65122 34700
rect 65613 34697 65625 34700
rect 65659 34697 65671 34731
rect 65613 34691 65671 34697
rect 66806 34688 66812 34740
rect 66864 34728 66870 34740
rect 67085 34731 67143 34737
rect 67085 34728 67097 34731
rect 66864 34700 67097 34728
rect 66864 34688 66870 34700
rect 67085 34697 67097 34700
rect 67131 34697 67143 34731
rect 67085 34691 67143 34697
rect 66349 34663 66407 34669
rect 66349 34629 66361 34663
rect 66395 34660 66407 34663
rect 67266 34660 67272 34672
rect 66395 34632 67272 34660
rect 66395 34629 66407 34632
rect 66349 34623 66407 34629
rect 67266 34620 67272 34632
rect 67324 34620 67330 34672
rect 63250 34536 63632 34564
rect 63604 34524 63632 34536
rect 65058 34524 65064 34536
rect 63604 34496 65064 34524
rect 65058 34484 65064 34496
rect 65116 34484 65122 34536
rect 66257 34527 66315 34533
rect 66257 34493 66269 34527
rect 66303 34524 66315 34527
rect 66346 34524 66352 34536
rect 66303 34496 66352 34524
rect 66303 34493 66315 34496
rect 66257 34487 66315 34493
rect 66346 34484 66352 34496
rect 66404 34484 66410 34536
rect 66806 34484 66812 34536
rect 66864 34524 66870 34536
rect 66901 34527 66959 34533
rect 66901 34524 66913 34527
rect 66864 34496 66913 34524
rect 66864 34484 66870 34496
rect 66901 34493 66913 34496
rect 66947 34493 66959 34527
rect 66901 34487 66959 34493
rect 67726 34484 67732 34536
rect 67784 34484 67790 34536
rect 65320 34298 74980 34320
rect 63236 33980 63264 34298
rect 65320 34246 71858 34298
rect 71910 34246 71922 34298
rect 71974 34246 71986 34298
rect 72038 34246 72050 34298
rect 72102 34246 72114 34298
rect 72166 34246 74980 34298
rect 65320 34224 74980 34246
rect 65613 34187 65671 34193
rect 65613 34153 65625 34187
rect 65659 34184 65671 34187
rect 65702 34184 65708 34196
rect 65659 34156 65708 34184
rect 65659 34153 65671 34156
rect 65613 34147 65671 34153
rect 65702 34144 65708 34156
rect 65760 34144 65766 34196
rect 66254 34144 66260 34196
rect 66312 34184 66318 34196
rect 66349 34187 66407 34193
rect 66349 34184 66361 34187
rect 66312 34156 66361 34184
rect 66312 34144 66318 34156
rect 66349 34153 66361 34156
rect 66395 34153 66407 34187
rect 66349 34147 66407 34153
rect 67085 34187 67143 34193
rect 67085 34153 67097 34187
rect 67131 34184 67143 34187
rect 67634 34184 67640 34196
rect 67131 34156 67640 34184
rect 67131 34153 67143 34156
rect 67085 34147 67143 34153
rect 67634 34144 67640 34156
rect 67692 34144 67698 34196
rect 66257 34051 66315 34057
rect 66257 34017 66269 34051
rect 66303 34048 66315 34051
rect 67082 34048 67088 34060
rect 66303 34020 67088 34048
rect 66303 34017 66315 34020
rect 66257 34011 66315 34017
rect 67082 34008 67088 34020
rect 67140 34008 67146 34060
rect 65150 33980 65156 33992
rect 63236 33952 65156 33980
rect 65150 33940 65156 33952
rect 65208 33940 65214 33992
rect 66990 33940 66996 33992
rect 67048 33940 67054 33992
rect 67729 33983 67787 33989
rect 67729 33949 67741 33983
rect 67775 33980 67787 33983
rect 68830 33980 68836 33992
rect 67775 33952 68836 33980
rect 67775 33949 67787 33952
rect 67729 33943 67787 33949
rect 68830 33940 68836 33952
rect 68888 33940 68894 33992
rect 65320 33754 74980 33776
rect 65320 33702 74210 33754
rect 74262 33702 74274 33754
rect 74326 33702 74338 33754
rect 74390 33702 74402 33754
rect 74454 33702 74466 33754
rect 74518 33702 74980 33754
rect 65320 33680 74980 33702
rect 65518 33600 65524 33652
rect 65576 33640 65582 33652
rect 65613 33643 65671 33649
rect 65613 33640 65625 33643
rect 65576 33612 65625 33640
rect 65576 33600 65582 33612
rect 65613 33609 65625 33612
rect 65659 33609 65671 33643
rect 65613 33603 65671 33609
rect 65702 33396 65708 33448
rect 65760 33436 65766 33448
rect 66165 33439 66223 33445
rect 66165 33436 66177 33439
rect 65760 33408 66177 33436
rect 65760 33396 65766 33408
rect 66165 33405 66177 33408
rect 66211 33405 66223 33439
rect 66165 33399 66223 33405
rect 63236 33300 63264 33322
rect 64874 33300 64880 33312
rect 63236 33272 64880 33300
rect 64874 33260 64880 33272
rect 64932 33260 64938 33312
rect 65320 33210 74980 33232
rect 65320 33158 71858 33210
rect 71910 33158 71922 33210
rect 71974 33158 71986 33210
rect 72038 33158 72050 33210
rect 72102 33158 72114 33210
rect 72166 33158 74980 33210
rect 65320 33136 74980 33158
rect 65613 33099 65671 33105
rect 65613 33065 65625 33099
rect 65659 33096 65671 33099
rect 66162 33096 66168 33108
rect 65659 33068 66168 33096
rect 65659 33065 65671 33068
rect 65613 33059 65671 33065
rect 66162 33056 66168 33068
rect 66220 33056 66226 33108
rect 66257 32895 66315 32901
rect 66257 32861 66269 32895
rect 66303 32892 66315 32895
rect 69290 32892 69296 32904
rect 66303 32864 69296 32892
rect 66303 32861 66315 32864
rect 66257 32855 66315 32861
rect 69290 32852 69296 32864
rect 69348 32852 69354 32904
rect 65320 32666 74980 32688
rect 65320 32614 74210 32666
rect 74262 32614 74274 32666
rect 74326 32614 74338 32666
rect 74390 32614 74402 32666
rect 74454 32614 74466 32666
rect 74518 32614 74980 32666
rect 65320 32592 74980 32614
rect 65613 32555 65671 32561
rect 65613 32521 65625 32555
rect 65659 32552 65671 32555
rect 69566 32552 69572 32564
rect 65659 32524 69572 32552
rect 65659 32521 65671 32524
rect 65613 32515 65671 32521
rect 69566 32512 69572 32524
rect 69624 32512 69630 32564
rect 63236 32212 63264 32370
rect 66257 32351 66315 32357
rect 66257 32317 66269 32351
rect 66303 32348 66315 32351
rect 70210 32348 70216 32360
rect 66303 32320 70216 32348
rect 66303 32317 66315 32320
rect 66257 32311 66315 32317
rect 70210 32308 70216 32320
rect 70268 32308 70274 32360
rect 65242 32212 65248 32224
rect 63236 32184 65248 32212
rect 65242 32172 65248 32184
rect 65300 32172 65306 32224
rect 65320 32122 74980 32144
rect 63236 31940 63264 32118
rect 65320 32070 71858 32122
rect 71910 32070 71922 32122
rect 71974 32070 71986 32122
rect 72038 32070 72050 32122
rect 72102 32070 72114 32122
rect 72166 32070 74980 32122
rect 65320 32048 74980 32070
rect 66257 32011 66315 32017
rect 66257 31977 66269 32011
rect 66303 32008 66315 32011
rect 69658 32008 69664 32020
rect 66303 31980 69664 32008
rect 66303 31977 66315 31980
rect 66257 31971 66315 31977
rect 69658 31968 69664 31980
rect 69716 31968 69722 32020
rect 67266 31940 67272 31952
rect 63236 31912 67272 31940
rect 67266 31900 67272 31912
rect 67324 31900 67330 31952
rect 65705 31807 65763 31813
rect 65705 31773 65717 31807
rect 65751 31804 65763 31807
rect 67818 31804 67824 31816
rect 65751 31776 67824 31804
rect 65751 31773 65763 31776
rect 65705 31767 65763 31773
rect 67818 31764 67824 31776
rect 67876 31764 67882 31816
rect 65320 31578 74980 31600
rect 65320 31526 74210 31578
rect 74262 31526 74274 31578
rect 74326 31526 74338 31578
rect 74390 31526 74402 31578
rect 74454 31526 74466 31578
rect 74518 31526 74980 31578
rect 65320 31504 74980 31526
rect 65334 31424 65340 31476
rect 65392 31464 65398 31476
rect 65613 31467 65671 31473
rect 65613 31464 65625 31467
rect 65392 31436 65625 31464
rect 65392 31424 65398 31436
rect 65613 31433 65625 31436
rect 65659 31433 65671 31467
rect 65613 31427 65671 31433
rect 66257 31263 66315 31269
rect 66257 31229 66269 31263
rect 66303 31260 66315 31263
rect 69382 31260 69388 31272
rect 66303 31232 69388 31260
rect 66303 31229 66315 31232
rect 66257 31223 66315 31229
rect 69382 31220 69388 31232
rect 69440 31220 69446 31272
rect 63236 31124 63264 31142
rect 64874 31124 64880 31136
rect 63236 31096 64880 31124
rect 64874 31084 64880 31096
rect 64932 31084 64938 31136
rect 65320 31034 74980 31056
rect 65320 30982 71858 31034
rect 71910 30982 71922 31034
rect 71974 30982 71986 31034
rect 72038 30982 72050 31034
rect 72102 30982 72114 31034
rect 72166 30982 74980 31034
rect 65320 30960 74980 30982
rect 66257 30923 66315 30929
rect 66257 30889 66269 30923
rect 66303 30920 66315 30923
rect 67174 30920 67180 30932
rect 66303 30892 67180 30920
rect 66303 30889 66315 30892
rect 66257 30883 66315 30889
rect 67174 30880 67180 30892
rect 67232 30880 67238 30932
rect 65705 30719 65763 30725
rect 65705 30685 65717 30719
rect 65751 30716 65763 30719
rect 69658 30716 69664 30728
rect 65751 30688 69664 30716
rect 65751 30685 65763 30688
rect 65705 30679 65763 30685
rect 69658 30676 69664 30688
rect 69716 30676 69722 30728
rect 65320 30490 74980 30512
rect 65320 30438 74210 30490
rect 74262 30438 74274 30490
rect 74326 30438 74338 30490
rect 74390 30438 74402 30490
rect 74454 30438 74466 30490
rect 74518 30438 74980 30490
rect 65320 30416 74980 30438
rect 65426 30268 65432 30320
rect 65484 30308 65490 30320
rect 65613 30311 65671 30317
rect 65613 30308 65625 30311
rect 65484 30280 65625 30308
rect 65484 30268 65490 30280
rect 65613 30277 65625 30280
rect 65659 30277 65671 30311
rect 65613 30271 65671 30277
rect 63236 30036 63264 30190
rect 66257 30175 66315 30181
rect 66257 30141 66269 30175
rect 66303 30172 66315 30175
rect 67174 30172 67180 30184
rect 66303 30144 67180 30172
rect 66303 30141 66315 30144
rect 66257 30135 66315 30141
rect 67174 30132 67180 30144
rect 67232 30132 67238 30184
rect 65334 30036 65340 30048
rect 63236 30008 65340 30036
rect 65334 29996 65340 30008
rect 65392 29996 65398 30048
rect 66254 29996 66260 30048
rect 66312 30036 66318 30048
rect 66714 30036 66720 30048
rect 66312 30008 66720 30036
rect 66312 29996 66318 30008
rect 66714 29996 66720 30008
rect 66772 29996 66778 30048
rect 65320 29946 74980 29968
rect 63236 29560 63264 29938
rect 65320 29894 71858 29946
rect 71910 29894 71922 29946
rect 71974 29894 71986 29946
rect 72038 29894 72050 29946
rect 72102 29894 72114 29946
rect 72166 29894 74980 29946
rect 65320 29872 74980 29894
rect 66257 29835 66315 29841
rect 66257 29801 66269 29835
rect 66303 29832 66315 29835
rect 66438 29832 66444 29844
rect 66303 29804 66444 29832
rect 66303 29801 66315 29804
rect 66257 29795 66315 29801
rect 66438 29792 66444 29804
rect 66496 29792 66502 29844
rect 65705 29631 65763 29637
rect 65705 29597 65717 29631
rect 65751 29628 65763 29631
rect 66162 29628 66168 29640
rect 65751 29600 66168 29628
rect 65751 29597 65763 29600
rect 65705 29591 65763 29597
rect 66162 29588 66168 29600
rect 66220 29588 66226 29640
rect 66438 29560 66444 29572
rect 63236 29532 66444 29560
rect 66438 29520 66444 29532
rect 66496 29520 66502 29572
rect 65320 29402 74980 29424
rect 65320 29350 74210 29402
rect 74262 29350 74274 29402
rect 74326 29350 74338 29402
rect 74390 29350 74402 29402
rect 74454 29350 74466 29402
rect 74518 29350 74980 29402
rect 65320 29328 74980 29350
rect 66254 29248 66260 29300
rect 66312 29248 66318 29300
rect 65705 29155 65763 29161
rect 65705 29121 65717 29155
rect 65751 29152 65763 29155
rect 69566 29152 69572 29164
rect 65751 29124 69572 29152
rect 65751 29121 65763 29124
rect 65705 29115 65763 29121
rect 69566 29112 69572 29124
rect 69624 29112 69630 29164
rect 66346 29044 66352 29096
rect 66404 29084 66410 29096
rect 67266 29084 67272 29096
rect 66404 29056 67272 29084
rect 66404 29044 66410 29056
rect 67266 29044 67272 29056
rect 67324 29044 67330 29096
rect 65150 28976 65156 29028
rect 65208 29016 65214 29028
rect 65208 28988 67312 29016
rect 65208 28976 65214 28988
rect 63236 28676 63264 28962
rect 67284 28960 67312 28988
rect 67266 28908 67272 28960
rect 67324 28908 67330 28960
rect 65320 28858 74980 28880
rect 65320 28806 71858 28858
rect 71910 28806 71922 28858
rect 71974 28806 71986 28858
rect 72038 28806 72050 28858
rect 72102 28806 72114 28858
rect 72166 28806 74980 28858
rect 65320 28784 74980 28806
rect 65610 28704 65616 28756
rect 65668 28744 65674 28756
rect 66901 28747 66959 28753
rect 66901 28744 66913 28747
rect 65668 28716 66913 28744
rect 65668 28704 65674 28716
rect 66901 28713 66913 28716
rect 66947 28744 66959 28747
rect 69106 28744 69112 28756
rect 66947 28716 69112 28744
rect 66947 28713 66959 28716
rect 66901 28707 66959 28713
rect 69106 28704 69112 28716
rect 69164 28704 69170 28756
rect 64874 28676 64880 28688
rect 63236 28648 64880 28676
rect 64874 28636 64880 28648
rect 64932 28636 64938 28688
rect 65613 28475 65671 28481
rect 65613 28441 65625 28475
rect 65659 28472 65671 28475
rect 66622 28472 66628 28484
rect 65659 28444 66628 28472
rect 65659 28441 65671 28444
rect 65613 28435 65671 28441
rect 66622 28432 66628 28444
rect 66680 28432 66686 28484
rect 65320 28314 74980 28336
rect 65320 28262 74210 28314
rect 74262 28262 74274 28314
rect 74326 28262 74338 28314
rect 74390 28262 74402 28314
rect 74454 28262 74466 28314
rect 74518 28262 74980 28314
rect 65320 28240 74980 28262
rect 65613 28203 65671 28209
rect 65613 28169 65625 28203
rect 65659 28200 65671 28203
rect 65978 28200 65984 28212
rect 65659 28172 65984 28200
rect 65659 28169 65671 28172
rect 65613 28163 65671 28169
rect 65978 28160 65984 28172
rect 66036 28160 66042 28212
rect 63236 27860 63264 28010
rect 66257 27999 66315 28005
rect 66257 27965 66269 27999
rect 66303 27996 66315 27999
rect 68002 27996 68008 28008
rect 66303 27968 68008 27996
rect 66303 27965 66315 27968
rect 66257 27959 66315 27965
rect 68002 27956 68008 27968
rect 68060 27956 68066 28008
rect 65518 27860 65524 27872
rect 63236 27832 65524 27860
rect 65518 27820 65524 27832
rect 65576 27820 65582 27872
rect 66622 27820 66628 27872
rect 66680 27860 66686 27872
rect 69014 27860 69020 27872
rect 66680 27832 69020 27860
rect 66680 27820 66686 27832
rect 69014 27820 69020 27832
rect 69072 27820 69078 27872
rect 65320 27770 74980 27792
rect 63236 27656 63264 27758
rect 65320 27718 71858 27770
rect 71910 27718 71922 27770
rect 71974 27718 71986 27770
rect 72038 27718 72050 27770
rect 72102 27718 72114 27770
rect 72166 27718 74980 27770
rect 65320 27696 74980 27718
rect 65150 27656 65156 27668
rect 63236 27628 65156 27656
rect 65150 27616 65156 27628
rect 65208 27616 65214 27668
rect 66349 27591 66407 27597
rect 66349 27557 66361 27591
rect 66395 27588 66407 27591
rect 66714 27588 66720 27600
rect 66395 27560 66720 27588
rect 66395 27557 66407 27560
rect 66349 27551 66407 27557
rect 66714 27548 66720 27560
rect 66772 27548 66778 27600
rect 64230 27480 64236 27532
rect 64288 27520 64294 27532
rect 66901 27523 66959 27529
rect 66901 27520 66913 27523
rect 64288 27492 66913 27520
rect 64288 27480 64294 27492
rect 66901 27489 66913 27492
rect 66947 27489 66959 27523
rect 66901 27483 66959 27489
rect 65794 27412 65800 27464
rect 65852 27452 65858 27464
rect 66257 27455 66315 27461
rect 66257 27452 66269 27455
rect 65852 27424 66269 27452
rect 65852 27412 65858 27424
rect 66257 27421 66269 27424
rect 66303 27421 66315 27455
rect 66257 27415 66315 27421
rect 65613 27387 65671 27393
rect 65613 27353 65625 27387
rect 65659 27384 65671 27387
rect 69750 27384 69756 27396
rect 65659 27356 69756 27384
rect 65659 27353 65671 27356
rect 65613 27347 65671 27353
rect 69750 27344 69756 27356
rect 69808 27344 69814 27396
rect 65320 27226 74980 27248
rect 65320 27174 74210 27226
rect 74262 27174 74274 27226
rect 74326 27174 74338 27226
rect 74390 27174 74402 27226
rect 74454 27174 74466 27226
rect 74518 27174 74980 27226
rect 65320 27152 74980 27174
rect 67085 27115 67143 27121
rect 67085 27081 67097 27115
rect 67131 27112 67143 27115
rect 67266 27112 67272 27124
rect 67131 27084 67272 27112
rect 67131 27081 67143 27084
rect 67085 27075 67143 27081
rect 67266 27072 67272 27084
rect 67324 27072 67330 27124
rect 66530 27004 66536 27056
rect 66588 27004 66594 27056
rect 64322 26936 64328 26988
rect 64380 26976 64386 26988
rect 65613 26979 65671 26985
rect 65613 26976 65625 26979
rect 64380 26948 65625 26976
rect 64380 26936 64386 26948
rect 65613 26945 65625 26948
rect 65659 26945 65671 26979
rect 65613 26939 65671 26945
rect 67729 26911 67787 26917
rect 67729 26877 67741 26911
rect 67775 26908 67787 26911
rect 68738 26908 68744 26920
rect 67775 26880 68744 26908
rect 67775 26877 67787 26880
rect 67729 26871 67787 26877
rect 68738 26868 68744 26880
rect 68796 26868 68802 26920
rect 63236 26772 63264 26782
rect 64874 26772 64880 26784
rect 63236 26744 64880 26772
rect 64874 26732 64880 26744
rect 64932 26772 64938 26784
rect 66438 26772 66444 26784
rect 64932 26744 66444 26772
rect 64932 26732 64938 26744
rect 66438 26732 66444 26744
rect 66496 26732 66502 26784
rect 65320 26682 74980 26704
rect 65320 26630 71858 26682
rect 71910 26630 71922 26682
rect 71974 26630 71986 26682
rect 72038 26630 72050 26682
rect 72102 26630 72114 26682
rect 72166 26630 74980 26682
rect 65320 26608 74980 26630
rect 65613 26571 65671 26577
rect 65613 26537 65625 26571
rect 65659 26568 65671 26571
rect 69198 26568 69204 26580
rect 65659 26540 69204 26568
rect 65659 26537 65671 26540
rect 65613 26531 65671 26537
rect 69198 26528 69204 26540
rect 69256 26528 69262 26580
rect 66257 26367 66315 26373
rect 66257 26333 66269 26367
rect 66303 26364 66315 26367
rect 67266 26364 67272 26376
rect 66303 26336 67272 26364
rect 66303 26333 66315 26336
rect 66257 26327 66315 26333
rect 67266 26324 67272 26336
rect 67324 26324 67330 26376
rect 65320 26138 74980 26160
rect 65320 26086 74210 26138
rect 74262 26086 74274 26138
rect 74326 26086 74338 26138
rect 74390 26086 74402 26138
rect 74454 26086 74466 26138
rect 74518 26086 74980 26138
rect 65320 26064 74980 26086
rect 65613 26027 65671 26033
rect 65613 25993 65625 26027
rect 65659 26024 65671 26027
rect 69842 26024 69848 26036
rect 65659 25996 69848 26024
rect 65659 25993 65671 25996
rect 65613 25987 65671 25993
rect 69842 25984 69848 25996
rect 69900 25984 69906 26036
rect 63236 25684 63264 25830
rect 66257 25823 66315 25829
rect 66257 25789 66269 25823
rect 66303 25820 66315 25823
rect 71498 25820 71504 25832
rect 66303 25792 71504 25820
rect 66303 25789 66315 25792
rect 66257 25783 66315 25789
rect 71498 25780 71504 25792
rect 71556 25780 71562 25832
rect 65426 25684 65432 25696
rect 63236 25656 65432 25684
rect 65426 25644 65432 25656
rect 65484 25644 65490 25696
rect 65320 25594 74980 25616
rect 63236 25276 63264 25578
rect 65320 25542 71858 25594
rect 71910 25542 71922 25594
rect 71974 25542 71986 25594
rect 72038 25542 72050 25594
rect 72102 25542 72114 25594
rect 72166 25542 74980 25594
rect 65320 25520 74980 25542
rect 65613 25483 65671 25489
rect 65613 25449 65625 25483
rect 65659 25480 65671 25483
rect 67450 25480 67456 25492
rect 65659 25452 67456 25480
rect 65659 25449 65671 25452
rect 65613 25443 65671 25449
rect 67450 25440 67456 25452
rect 67508 25440 67514 25492
rect 67082 25372 67088 25424
rect 67140 25412 67146 25424
rect 67140 25384 67496 25412
rect 67140 25372 67146 25384
rect 67468 25356 67496 25384
rect 67450 25304 67456 25356
rect 67508 25304 67514 25356
rect 65978 25276 65984 25288
rect 63236 25248 65984 25276
rect 65978 25236 65984 25248
rect 66036 25236 66042 25288
rect 66257 25279 66315 25285
rect 66257 25245 66269 25279
rect 66303 25276 66315 25279
rect 67082 25276 67088 25288
rect 66303 25248 67088 25276
rect 66303 25245 66315 25248
rect 66257 25239 66315 25245
rect 67082 25236 67088 25248
rect 67140 25236 67146 25288
rect 65320 25050 74980 25072
rect 65320 24998 74210 25050
rect 74262 24998 74274 25050
rect 74326 24998 74338 25050
rect 74390 24998 74402 25050
rect 74454 24998 74466 25050
rect 74518 24998 74980 25050
rect 65320 24976 74980 24998
rect 65610 24828 65616 24880
rect 65668 24868 65674 24880
rect 66254 24868 66260 24880
rect 65668 24840 66260 24868
rect 65668 24828 65674 24840
rect 66254 24828 66260 24840
rect 66312 24828 66318 24880
rect 66346 24760 66352 24812
rect 66404 24760 66410 24812
rect 66254 24692 66260 24744
rect 66312 24692 66318 24744
rect 66993 24735 67051 24741
rect 66993 24701 67005 24735
rect 67039 24732 67051 24735
rect 69750 24732 69756 24744
rect 67039 24704 69756 24732
rect 67039 24701 67051 24704
rect 66993 24695 67051 24701
rect 69750 24692 69756 24704
rect 69808 24692 69814 24744
rect 65613 24667 65671 24673
rect 65613 24633 65625 24667
rect 65659 24664 65671 24667
rect 67358 24664 67364 24676
rect 65659 24636 67364 24664
rect 65659 24633 65671 24636
rect 65613 24627 65671 24633
rect 67358 24624 67364 24636
rect 67416 24624 67422 24676
rect 63236 24324 63264 24602
rect 65320 24506 74980 24528
rect 65320 24454 71858 24506
rect 71910 24454 71922 24506
rect 71974 24454 71986 24506
rect 72038 24454 72050 24506
rect 72102 24454 72114 24506
rect 72166 24454 74980 24506
rect 65320 24432 74980 24454
rect 65613 24395 65671 24401
rect 65613 24361 65625 24395
rect 65659 24392 65671 24395
rect 66898 24392 66904 24404
rect 65659 24364 66904 24392
rect 65659 24361 65671 24364
rect 65613 24355 65671 24361
rect 66898 24352 66904 24364
rect 66956 24352 66962 24404
rect 66993 24395 67051 24401
rect 66993 24361 67005 24395
rect 67039 24392 67051 24395
rect 68370 24392 68376 24404
rect 67039 24364 68376 24392
rect 67039 24361 67051 24364
rect 66993 24355 67051 24361
rect 68370 24352 68376 24364
rect 68428 24352 68434 24404
rect 64874 24324 64880 24336
rect 63236 24296 64880 24324
rect 64874 24284 64880 24296
rect 64932 24284 64938 24336
rect 66257 24259 66315 24265
rect 66257 24225 66269 24259
rect 66303 24256 66315 24259
rect 66530 24256 66536 24268
rect 66303 24228 66536 24256
rect 66303 24225 66315 24228
rect 66257 24219 66315 24225
rect 66530 24216 66536 24228
rect 66588 24216 66594 24268
rect 66346 24148 66352 24200
rect 66404 24148 66410 24200
rect 65320 23962 74980 23984
rect 65320 23910 74210 23962
rect 74262 23910 74274 23962
rect 74326 23910 74338 23962
rect 74390 23910 74402 23962
rect 74454 23910 74466 23962
rect 74518 23910 74980 23962
rect 65320 23888 74980 23910
rect 65610 23808 65616 23860
rect 65668 23808 65674 23860
rect 66349 23851 66407 23857
rect 66349 23817 66361 23851
rect 66395 23848 66407 23851
rect 66806 23848 66812 23860
rect 66395 23820 66812 23848
rect 66395 23817 66407 23820
rect 66349 23811 66407 23817
rect 66806 23808 66812 23820
rect 66864 23808 66870 23860
rect 67085 23851 67143 23857
rect 67085 23817 67097 23851
rect 67131 23848 67143 23851
rect 67726 23848 67732 23860
rect 67131 23820 67732 23848
rect 67131 23817 67143 23820
rect 67085 23811 67143 23817
rect 67726 23808 67732 23820
rect 67784 23808 67790 23860
rect 64874 23672 64880 23724
rect 64932 23712 64938 23724
rect 65610 23712 65616 23724
rect 64932 23684 65616 23712
rect 64932 23672 64938 23684
rect 65610 23672 65616 23684
rect 65668 23672 65674 23724
rect 63236 23508 63264 23650
rect 66257 23647 66315 23653
rect 66257 23613 66269 23647
rect 66303 23644 66315 23647
rect 66622 23644 66628 23656
rect 66303 23616 66628 23644
rect 66303 23613 66315 23616
rect 66257 23607 66315 23613
rect 66622 23604 66628 23616
rect 66680 23604 66686 23656
rect 66806 23604 66812 23656
rect 66864 23644 66870 23656
rect 66901 23647 66959 23653
rect 66901 23644 66913 23647
rect 66864 23616 66913 23644
rect 66864 23604 66870 23616
rect 66901 23613 66913 23616
rect 66947 23613 66959 23647
rect 66901 23607 66959 23613
rect 67729 23647 67787 23653
rect 67729 23613 67741 23647
rect 67775 23644 67787 23647
rect 68922 23644 68928 23656
rect 67775 23616 68928 23644
rect 67775 23613 67787 23616
rect 67729 23607 67787 23613
rect 68922 23604 68928 23616
rect 68980 23604 68986 23656
rect 64874 23508 64880 23520
rect 63236 23480 64880 23508
rect 64874 23468 64880 23480
rect 64932 23468 64938 23520
rect 65320 23418 74980 23440
rect 63236 23032 63264 23398
rect 65320 23366 71858 23418
rect 71910 23366 71922 23418
rect 71974 23366 71986 23418
rect 72038 23366 72050 23418
rect 72102 23366 72114 23418
rect 72166 23366 74980 23418
rect 65320 23344 74980 23366
rect 66714 23264 66720 23316
rect 66772 23304 66778 23316
rect 67085 23307 67143 23313
rect 67085 23304 67097 23307
rect 66772 23276 67097 23304
rect 66772 23264 66778 23276
rect 67085 23273 67097 23276
rect 67131 23273 67143 23307
rect 67085 23267 67143 23273
rect 66349 23239 66407 23245
rect 66349 23205 66361 23239
rect 66395 23236 66407 23239
rect 66990 23236 66996 23248
rect 66395 23208 66996 23236
rect 66395 23205 66407 23208
rect 66349 23199 66407 23205
rect 66990 23196 66996 23208
rect 67048 23196 67054 23248
rect 66257 23171 66315 23177
rect 66257 23137 66269 23171
rect 66303 23168 66315 23171
rect 67358 23168 67364 23180
rect 66303 23140 67364 23168
rect 66303 23137 66315 23140
rect 66257 23131 66315 23137
rect 67358 23128 67364 23140
rect 67416 23128 67422 23180
rect 66898 23060 66904 23112
rect 66956 23060 66962 23112
rect 67729 23103 67787 23109
rect 67729 23069 67741 23103
rect 67775 23100 67787 23103
rect 67910 23100 67916 23112
rect 67775 23072 67916 23100
rect 67775 23069 67787 23072
rect 67729 23063 67787 23069
rect 67910 23060 67916 23072
rect 67968 23060 67974 23112
rect 65426 23032 65432 23044
rect 63236 23004 65432 23032
rect 65426 22992 65432 23004
rect 65484 22992 65490 23044
rect 65613 23035 65671 23041
rect 65613 23001 65625 23035
rect 65659 23032 65671 23035
rect 67450 23032 67456 23044
rect 65659 23004 67456 23032
rect 65659 23001 65671 23004
rect 65613 22995 65671 23001
rect 67450 22992 67456 23004
rect 67508 22992 67514 23044
rect 65320 22874 74980 22896
rect 65320 22822 74210 22874
rect 74262 22822 74274 22874
rect 74326 22822 74338 22874
rect 74390 22822 74402 22874
rect 74454 22822 74466 22874
rect 74518 22822 74980 22874
rect 65320 22800 74980 22822
rect 65613 22763 65671 22769
rect 65613 22729 65625 22763
rect 65659 22760 65671 22763
rect 65702 22760 65708 22772
rect 65659 22732 65708 22760
rect 65659 22729 65671 22732
rect 65613 22723 65671 22729
rect 65702 22720 65708 22732
rect 65760 22720 65766 22772
rect 66257 22559 66315 22565
rect 66257 22525 66269 22559
rect 66303 22556 66315 22559
rect 66714 22556 66720 22568
rect 66303 22528 66720 22556
rect 66303 22525 66315 22528
rect 66257 22519 66315 22525
rect 66714 22516 66720 22528
rect 66772 22516 66778 22568
rect 63236 22148 63264 22422
rect 65320 22330 74980 22352
rect 65320 22278 71858 22330
rect 71910 22278 71922 22330
rect 71974 22278 71986 22330
rect 72038 22278 72050 22330
rect 72102 22278 72114 22330
rect 72166 22278 74980 22330
rect 65320 22256 74980 22278
rect 65702 22148 65708 22160
rect 63236 22120 65708 22148
rect 65702 22108 65708 22120
rect 65760 22108 65766 22160
rect 66438 22040 66444 22092
rect 66496 22040 66502 22092
rect 68554 22040 68560 22092
rect 68612 22080 68618 22092
rect 68649 22083 68707 22089
rect 68649 22080 68661 22083
rect 68612 22052 68661 22080
rect 68612 22040 68618 22052
rect 68649 22049 68661 22052
rect 68695 22049 68707 22083
rect 68649 22043 68707 22049
rect 70118 22040 70124 22092
rect 70176 22040 70182 22092
rect 65797 22015 65855 22021
rect 65797 21981 65809 22015
rect 65843 22012 65855 22015
rect 67634 22012 67640 22024
rect 65843 21984 67640 22012
rect 65843 21981 65855 21984
rect 65797 21975 65855 21981
rect 67634 21972 67640 21984
rect 67692 21972 67698 22024
rect 69293 22015 69351 22021
rect 69293 21981 69305 22015
rect 69339 22012 69351 22015
rect 69934 22012 69940 22024
rect 69339 21984 69940 22012
rect 69339 21981 69351 21984
rect 69293 21975 69351 21981
rect 69934 21972 69940 21984
rect 69992 21972 69998 22024
rect 70765 22015 70823 22021
rect 70765 21981 70777 22015
rect 70811 22012 70823 22015
rect 71590 22012 71596 22024
rect 70811 21984 71596 22012
rect 70811 21981 70823 21984
rect 70765 21975 70823 21981
rect 71590 21972 71596 21984
rect 71648 21972 71654 22024
rect 65320 21786 74980 21808
rect 65320 21734 74210 21786
rect 74262 21734 74274 21786
rect 74326 21734 74338 21786
rect 74390 21734 74402 21786
rect 74454 21734 74466 21786
rect 74518 21734 74980 21786
rect 65320 21712 74980 21734
rect 65150 21632 65156 21684
rect 65208 21672 65214 21684
rect 65613 21675 65671 21681
rect 65613 21672 65625 21675
rect 65208 21644 65625 21672
rect 65208 21632 65214 21644
rect 65613 21641 65625 21644
rect 65659 21641 65671 21675
rect 65613 21635 65671 21641
rect 66257 21471 66315 21477
rect 63236 21332 63264 21470
rect 66257 21437 66269 21471
rect 66303 21468 66315 21471
rect 69842 21468 69848 21480
rect 66303 21440 69848 21468
rect 66303 21437 66315 21440
rect 66257 21431 66315 21437
rect 69842 21428 69848 21440
rect 69900 21428 69906 21480
rect 65150 21360 65156 21412
rect 65208 21400 65214 21412
rect 65518 21400 65524 21412
rect 65208 21372 65524 21400
rect 65208 21360 65214 21372
rect 65518 21360 65524 21372
rect 65576 21360 65582 21412
rect 64782 21332 64788 21344
rect 63236 21304 64788 21332
rect 64782 21292 64788 21304
rect 64840 21292 64846 21344
rect 65320 21242 74980 21264
rect 63236 20924 63264 21218
rect 65320 21190 71858 21242
rect 71910 21190 71922 21242
rect 71974 21190 71986 21242
rect 72038 21190 72050 21242
rect 72102 21190 72114 21242
rect 72166 21190 74980 21242
rect 65320 21168 74980 21190
rect 68186 21088 68192 21140
rect 68244 21088 68250 21140
rect 65610 20924 65616 20936
rect 63236 20896 65616 20924
rect 65610 20884 65616 20896
rect 65668 20884 65674 20936
rect 68833 20927 68891 20933
rect 68833 20893 68845 20927
rect 68879 20924 68891 20927
rect 70118 20924 70124 20936
rect 68879 20896 70124 20924
rect 68879 20893 68891 20896
rect 68833 20887 68891 20893
rect 70118 20884 70124 20896
rect 70176 20884 70182 20936
rect 66254 20748 66260 20800
rect 66312 20788 66318 20800
rect 67450 20788 67456 20800
rect 66312 20760 67456 20788
rect 66312 20748 66318 20760
rect 67450 20748 67456 20760
rect 67508 20748 67514 20800
rect 65320 20698 74980 20720
rect 65320 20646 74210 20698
rect 74262 20646 74274 20698
rect 74326 20646 74338 20698
rect 74390 20646 74402 20698
rect 74454 20646 74466 20698
rect 74518 20646 74980 20698
rect 65320 20624 74980 20646
rect 67085 20587 67143 20593
rect 67085 20553 67097 20587
rect 67131 20584 67143 20587
rect 67542 20584 67548 20596
rect 67131 20556 67548 20584
rect 67131 20553 67143 20556
rect 67085 20547 67143 20553
rect 67542 20544 67548 20556
rect 67600 20544 67606 20596
rect 66349 20519 66407 20525
rect 66349 20485 66361 20519
rect 66395 20516 66407 20519
rect 69474 20516 69480 20528
rect 66395 20488 69480 20516
rect 66395 20485 66407 20488
rect 66349 20479 66407 20485
rect 69474 20476 69480 20488
rect 69532 20476 69538 20528
rect 66993 20451 67051 20457
rect 66993 20417 67005 20451
rect 67039 20448 67051 20451
rect 68278 20448 68284 20460
rect 67039 20420 68284 20448
rect 67039 20417 67051 20420
rect 66993 20411 67051 20417
rect 68278 20408 68284 20420
rect 68336 20408 68342 20460
rect 66257 20383 66315 20389
rect 66257 20349 66269 20383
rect 66303 20380 66315 20383
rect 67729 20383 67787 20389
rect 66303 20352 67036 20380
rect 66303 20349 66315 20352
rect 66257 20343 66315 20349
rect 67008 20324 67036 20352
rect 67729 20349 67741 20383
rect 67775 20380 67787 20383
rect 68370 20380 68376 20392
rect 67775 20352 68376 20380
rect 67775 20349 67787 20352
rect 67729 20343 67787 20349
rect 68370 20340 68376 20352
rect 68428 20340 68434 20392
rect 65702 20312 65708 20324
rect 64846 20284 65708 20312
rect 64846 20244 64874 20284
rect 65702 20272 65708 20284
rect 65760 20272 65766 20324
rect 66990 20272 66996 20324
rect 67048 20272 67054 20324
rect 63236 20216 64874 20244
rect 65613 20247 65671 20253
rect 65613 20213 65625 20247
rect 65659 20244 65671 20247
rect 70026 20244 70032 20256
rect 65659 20216 70032 20244
rect 65659 20213 65671 20216
rect 65613 20207 65671 20213
rect 70026 20204 70032 20216
rect 70084 20204 70090 20256
rect 65320 20154 74980 20176
rect 65320 20102 71858 20154
rect 71910 20102 71922 20154
rect 71974 20102 71986 20154
rect 72038 20102 72050 20154
rect 72102 20102 72114 20154
rect 72166 20102 74980 20154
rect 65320 20080 74980 20102
rect 65613 20043 65671 20049
rect 65613 20009 65625 20043
rect 65659 20040 65671 20043
rect 65978 20040 65984 20052
rect 65659 20012 65984 20040
rect 65659 20009 65671 20012
rect 65613 20003 65671 20009
rect 65978 20000 65984 20012
rect 66036 20000 66042 20052
rect 66622 19932 66628 19984
rect 66680 19972 66686 19984
rect 67082 19972 67088 19984
rect 66680 19944 67088 19972
rect 66680 19932 66686 19944
rect 67082 19932 67088 19944
rect 67140 19932 67146 19984
rect 65518 19864 65524 19916
rect 65576 19904 65582 19916
rect 65978 19904 65984 19916
rect 65576 19876 65984 19904
rect 65576 19864 65582 19876
rect 65978 19864 65984 19876
rect 66036 19864 66042 19916
rect 66257 19839 66315 19845
rect 66257 19805 66269 19839
rect 66303 19836 66315 19839
rect 69474 19836 69480 19848
rect 66303 19808 69480 19836
rect 66303 19805 66315 19808
rect 66257 19799 66315 19805
rect 69474 19796 69480 19808
rect 69532 19796 69538 19848
rect 65320 19610 74980 19632
rect 65320 19558 74210 19610
rect 74262 19558 74274 19610
rect 74326 19558 74338 19610
rect 74390 19558 74402 19610
rect 74454 19558 74466 19610
rect 74518 19558 74980 19610
rect 65320 19536 74980 19558
rect 66257 19499 66315 19505
rect 66257 19465 66269 19499
rect 66303 19496 66315 19499
rect 68186 19496 68192 19508
rect 66303 19468 68192 19496
rect 66303 19465 66315 19468
rect 66257 19459 66315 19465
rect 68186 19456 68192 19468
rect 68244 19456 68250 19508
rect 65705 19295 65763 19301
rect 63236 19224 63264 19290
rect 65705 19261 65717 19295
rect 65751 19292 65763 19295
rect 68554 19292 68560 19304
rect 65751 19264 68560 19292
rect 65751 19261 65763 19264
rect 65705 19255 65763 19261
rect 68554 19252 68560 19264
rect 68612 19252 68618 19304
rect 72326 19224 72332 19236
rect 63236 19196 72332 19224
rect 72326 19184 72332 19196
rect 72384 19184 72390 19236
rect 65320 19066 74980 19088
rect 63236 18748 63264 19038
rect 65320 19014 71858 19066
rect 71910 19014 71922 19066
rect 71974 19014 71986 19066
rect 72038 19014 72050 19066
rect 72102 19014 72114 19066
rect 72166 19014 74980 19066
rect 65320 18992 74980 19014
rect 66257 18955 66315 18961
rect 66257 18921 66269 18955
rect 66303 18952 66315 18955
rect 68462 18952 68468 18964
rect 66303 18924 68468 18952
rect 66303 18921 66315 18924
rect 66257 18915 66315 18921
rect 68462 18912 68468 18924
rect 68520 18912 68526 18964
rect 65518 18748 65524 18760
rect 63236 18720 65524 18748
rect 65518 18708 65524 18720
rect 65576 18708 65582 18760
rect 65705 18751 65763 18757
rect 65705 18717 65717 18751
rect 65751 18748 65763 18751
rect 72418 18748 72424 18760
rect 65751 18720 72424 18748
rect 65751 18717 65763 18720
rect 65705 18711 65763 18717
rect 72418 18708 72424 18720
rect 72476 18708 72482 18760
rect 65320 18522 74980 18544
rect 65320 18470 74210 18522
rect 74262 18470 74274 18522
rect 74326 18470 74338 18522
rect 74390 18470 74402 18522
rect 74454 18470 74466 18522
rect 74518 18470 74980 18522
rect 65320 18448 74980 18470
rect 65426 18368 65432 18420
rect 65484 18408 65490 18420
rect 65613 18411 65671 18417
rect 65613 18408 65625 18411
rect 65484 18380 65625 18408
rect 65484 18368 65490 18380
rect 65613 18377 65625 18380
rect 65659 18377 65671 18411
rect 65613 18371 65671 18377
rect 64874 18232 64880 18284
rect 64932 18272 64938 18284
rect 65426 18272 65432 18284
rect 64932 18244 65432 18272
rect 64932 18232 64938 18244
rect 65426 18232 65432 18244
rect 65484 18232 65490 18284
rect 66257 18207 66315 18213
rect 66257 18173 66269 18207
rect 66303 18204 66315 18207
rect 69198 18204 69204 18216
rect 66303 18176 69204 18204
rect 66303 18173 66315 18176
rect 66257 18167 66315 18173
rect 69198 18164 69204 18176
rect 69256 18164 69262 18216
rect 65702 18068 65708 18080
rect 63236 18040 65708 18068
rect 65702 18028 65708 18040
rect 65760 18028 65766 18080
rect 65320 17978 74980 18000
rect 65320 17926 71858 17978
rect 71910 17926 71922 17978
rect 71974 17926 71986 17978
rect 72038 17926 72050 17978
rect 72102 17926 72114 17978
rect 72166 17926 74980 17978
rect 65320 17904 74980 17926
rect 66257 17867 66315 17873
rect 66257 17833 66269 17867
rect 66303 17864 66315 17867
rect 68830 17864 68836 17876
rect 66303 17836 68836 17864
rect 66303 17833 66315 17836
rect 66257 17827 66315 17833
rect 68830 17824 68836 17836
rect 68888 17824 68894 17876
rect 65705 17663 65763 17669
rect 65705 17629 65717 17663
rect 65751 17660 65763 17663
rect 70578 17660 70584 17672
rect 65751 17632 70584 17660
rect 65751 17629 65763 17632
rect 65705 17623 65763 17629
rect 70578 17620 70584 17632
rect 70636 17620 70642 17672
rect 65320 17434 74980 17456
rect 65320 17382 74210 17434
rect 74262 17382 74274 17434
rect 74326 17382 74338 17434
rect 74390 17382 74402 17434
rect 74454 17382 74466 17434
rect 74518 17382 74980 17434
rect 65320 17360 74980 17382
rect 65610 17280 65616 17332
rect 65668 17280 65674 17332
rect 66349 17323 66407 17329
rect 66349 17289 66361 17323
rect 66395 17320 66407 17323
rect 70210 17320 70216 17332
rect 66395 17292 70216 17320
rect 66395 17289 66407 17292
rect 66349 17283 66407 17289
rect 70210 17280 70216 17292
rect 70268 17280 70274 17332
rect 70486 17184 70492 17196
rect 63604 17156 70492 17184
rect 63604 17124 63632 17156
rect 70486 17144 70492 17156
rect 70544 17144 70550 17196
rect 63250 17096 63632 17124
rect 66254 17076 66260 17128
rect 66312 17076 66318 17128
rect 66993 17119 67051 17125
rect 66993 17085 67005 17119
rect 67039 17116 67051 17119
rect 72234 17116 72240 17128
rect 67039 17088 72240 17116
rect 67039 17085 67051 17088
rect 66993 17079 67051 17085
rect 72234 17076 72240 17088
rect 72292 17076 72298 17128
rect 65320 16890 74980 16912
rect 63236 16640 63264 16858
rect 65320 16838 71858 16890
rect 71910 16838 71922 16890
rect 71974 16838 71986 16890
rect 72038 16838 72050 16890
rect 72102 16838 72114 16890
rect 72166 16838 74980 16890
rect 65320 16816 74980 16838
rect 64874 16640 64880 16652
rect 63236 16612 64880 16640
rect 64874 16600 64880 16612
rect 64932 16600 64938 16652
rect 66257 16643 66315 16649
rect 66257 16609 66269 16643
rect 66303 16640 66315 16643
rect 72510 16640 72516 16652
rect 66303 16612 72516 16640
rect 66303 16609 66315 16612
rect 66257 16603 66315 16609
rect 72510 16600 72516 16612
rect 72568 16600 72574 16652
rect 65613 16575 65671 16581
rect 65613 16541 65625 16575
rect 65659 16572 65671 16575
rect 67818 16572 67824 16584
rect 65659 16544 67824 16572
rect 65659 16541 65671 16544
rect 65613 16535 65671 16541
rect 67818 16532 67824 16544
rect 67876 16532 67882 16584
rect 65320 16346 74980 16368
rect 65320 16294 74210 16346
rect 74262 16294 74274 16346
rect 74326 16294 74338 16346
rect 74390 16294 74402 16346
rect 74454 16294 74466 16346
rect 74518 16294 74980 16346
rect 65320 16272 74980 16294
rect 65613 16235 65671 16241
rect 65613 16201 65625 16235
rect 65659 16232 65671 16235
rect 66162 16232 66168 16244
rect 65659 16204 66168 16232
rect 65659 16201 65671 16204
rect 65613 16195 65671 16201
rect 66162 16192 66168 16204
rect 66220 16192 66226 16244
rect 64690 16056 64696 16108
rect 64748 16096 64754 16108
rect 66990 16096 66996 16108
rect 64748 16068 66996 16096
rect 64748 16056 64754 16068
rect 66990 16056 66996 16068
rect 67048 16056 67054 16108
rect 66257 16031 66315 16037
rect 66257 15997 66269 16031
rect 66303 16028 66315 16031
rect 70394 16028 70400 16040
rect 66303 16000 70400 16028
rect 66303 15997 66315 16000
rect 66257 15991 66315 15997
rect 70394 15988 70400 16000
rect 70452 15988 70458 16040
rect 63236 15620 63264 15882
rect 65320 15802 74980 15824
rect 65320 15750 71858 15802
rect 71910 15750 71922 15802
rect 71974 15750 71986 15802
rect 72038 15750 72050 15802
rect 72102 15750 72114 15802
rect 72166 15750 74980 15802
rect 65320 15728 74980 15750
rect 65613 15691 65671 15697
rect 65613 15657 65625 15691
rect 65659 15688 65671 15691
rect 69658 15688 69664 15700
rect 65659 15660 69664 15688
rect 65659 15657 65671 15660
rect 65613 15651 65671 15657
rect 69658 15648 69664 15660
rect 69716 15648 69722 15700
rect 63236 15592 64874 15620
rect 64846 15552 64874 15592
rect 65610 15552 65616 15564
rect 64846 15524 65616 15552
rect 65610 15512 65616 15524
rect 65668 15512 65674 15564
rect 66257 15487 66315 15493
rect 66257 15453 66269 15487
rect 66303 15484 66315 15487
rect 70946 15484 70952 15496
rect 66303 15456 70952 15484
rect 66303 15453 66315 15456
rect 66257 15447 66315 15453
rect 70946 15444 70952 15456
rect 71004 15444 71010 15496
rect 65702 15308 65708 15360
rect 65760 15348 65766 15360
rect 66254 15348 66260 15360
rect 65760 15320 66260 15348
rect 65760 15308 65766 15320
rect 66254 15308 66260 15320
rect 66312 15308 66318 15360
rect 67542 15308 67548 15360
rect 67600 15348 67606 15360
rect 70762 15348 70768 15360
rect 67600 15320 70768 15348
rect 67600 15308 67606 15320
rect 70762 15308 70768 15320
rect 70820 15308 70826 15360
rect 65320 15258 74980 15280
rect 65320 15206 74210 15258
rect 74262 15206 74274 15258
rect 74326 15206 74338 15258
rect 74390 15206 74402 15258
rect 74454 15206 74466 15258
rect 74518 15206 74980 15258
rect 65320 15184 74980 15206
rect 65613 15147 65671 15153
rect 65613 15113 65625 15147
rect 65659 15144 65671 15147
rect 69566 15144 69572 15156
rect 65659 15116 69572 15144
rect 65659 15113 65671 15116
rect 65613 15107 65671 15113
rect 69566 15104 69572 15116
rect 69624 15104 69630 15156
rect 66257 14943 66315 14949
rect 63236 14912 64874 14940
rect 64846 14872 64874 14912
rect 66257 14909 66269 14943
rect 66303 14940 66315 14943
rect 69658 14940 69664 14952
rect 66303 14912 69664 14940
rect 66303 14909 66315 14912
rect 66257 14903 66315 14909
rect 69658 14900 69664 14912
rect 69716 14900 69722 14952
rect 72602 14872 72608 14884
rect 64846 14844 72608 14872
rect 72602 14832 72608 14844
rect 72660 14832 72666 14884
rect 65320 14714 74980 14736
rect 63236 14396 63264 14678
rect 65320 14662 71858 14714
rect 71910 14662 71922 14714
rect 71974 14662 71986 14714
rect 72038 14662 72050 14714
rect 72102 14662 72114 14714
rect 72166 14662 74980 14714
rect 65320 14640 74980 14662
rect 65518 14560 65524 14612
rect 65576 14600 65582 14612
rect 65613 14603 65671 14609
rect 65613 14600 65625 14603
rect 65576 14572 65625 14600
rect 65576 14560 65582 14572
rect 65613 14569 65625 14572
rect 65659 14569 65671 14603
rect 65613 14563 65671 14569
rect 69382 14492 69388 14544
rect 69440 14532 69446 14544
rect 69566 14532 69572 14544
rect 69440 14504 69572 14532
rect 69440 14492 69446 14504
rect 69566 14492 69572 14504
rect 69624 14492 69630 14544
rect 65610 14396 65616 14408
rect 63236 14368 65616 14396
rect 65610 14356 65616 14368
rect 65668 14356 65674 14408
rect 66257 14399 66315 14405
rect 66257 14365 66269 14399
rect 66303 14396 66315 14399
rect 67726 14396 67732 14408
rect 66303 14368 67732 14396
rect 66303 14365 66315 14368
rect 66257 14359 66315 14365
rect 67726 14356 67732 14368
rect 67784 14356 67790 14408
rect 65320 14170 74980 14192
rect 65320 14118 74210 14170
rect 74262 14118 74274 14170
rect 74326 14118 74338 14170
rect 74390 14118 74402 14170
rect 74454 14118 74466 14170
rect 74518 14118 74980 14170
rect 65320 14096 74980 14118
rect 63236 13376 63264 13702
rect 65320 13626 74980 13648
rect 65320 13574 71858 13626
rect 71910 13574 71922 13626
rect 71974 13574 71986 13626
rect 72038 13574 72050 13626
rect 72102 13574 72114 13626
rect 72166 13574 74980 13626
rect 65320 13552 74980 13574
rect 64874 13472 64880 13524
rect 64932 13512 64938 13524
rect 65613 13515 65671 13521
rect 65613 13512 65625 13515
rect 64932 13484 65625 13512
rect 64932 13472 64938 13484
rect 65613 13481 65625 13484
rect 65659 13481 65671 13515
rect 65613 13475 65671 13481
rect 64874 13376 64880 13388
rect 63236 13348 64880 13376
rect 64874 13336 64880 13348
rect 64932 13376 64938 13388
rect 65518 13376 65524 13388
rect 64932 13348 65524 13376
rect 64932 13336 64938 13348
rect 65518 13336 65524 13348
rect 65576 13336 65582 13388
rect 66257 13311 66315 13317
rect 66257 13277 66269 13311
rect 66303 13308 66315 13311
rect 68094 13308 68100 13320
rect 66303 13280 68100 13308
rect 66303 13277 66315 13280
rect 66257 13271 66315 13277
rect 68094 13268 68100 13280
rect 68152 13268 68158 13320
rect 65320 13082 74980 13104
rect 65320 13030 74210 13082
rect 74262 13030 74274 13082
rect 74326 13030 74338 13082
rect 74390 13030 74402 13082
rect 74454 13030 74466 13082
rect 74518 13030 74980 13082
rect 65320 13008 74980 13030
rect 65518 12764 65524 12776
rect 63250 12736 65524 12764
rect 65518 12724 65524 12736
rect 65576 12724 65582 12776
rect 66162 12628 66168 12640
rect 63236 12600 66168 12628
rect 63236 12498 63264 12600
rect 66162 12588 66168 12600
rect 66220 12588 66226 12640
rect 65320 12538 74980 12560
rect 65320 12486 71858 12538
rect 71910 12486 71922 12538
rect 71974 12486 71986 12538
rect 72038 12486 72050 12538
rect 72102 12486 72114 12538
rect 72166 12486 74980 12538
rect 65320 12464 74980 12486
rect 65320 11994 74980 12016
rect 65320 11942 74210 11994
rect 74262 11942 74274 11994
rect 74326 11942 74338 11994
rect 74390 11942 74402 11994
rect 74454 11942 74466 11994
rect 74518 11942 74980 11994
rect 65320 11920 74980 11942
rect 65610 11840 65616 11892
rect 65668 11840 65674 11892
rect 66257 11679 66315 11685
rect 66257 11645 66269 11679
rect 66303 11676 66315 11679
rect 69198 11676 69204 11688
rect 66303 11648 69204 11676
rect 66303 11645 66315 11648
rect 66257 11639 66315 11645
rect 69198 11636 69204 11648
rect 69256 11636 69262 11688
rect 63236 11268 63264 11522
rect 64966 11500 64972 11552
rect 65024 11540 65030 11552
rect 65518 11540 65524 11552
rect 65024 11512 65524 11540
rect 65024 11500 65030 11512
rect 65518 11500 65524 11512
rect 65576 11500 65582 11552
rect 63862 11432 63868 11484
rect 63920 11472 63926 11484
rect 64506 11472 64512 11484
rect 63920 11444 64512 11472
rect 63920 11432 63926 11444
rect 64506 11432 64512 11444
rect 64564 11432 64570 11484
rect 65320 11450 74980 11472
rect 63494 11364 63500 11416
rect 63552 11404 63558 11416
rect 64322 11404 64328 11416
rect 63552 11376 64328 11404
rect 63552 11364 63558 11376
rect 64322 11364 64328 11376
rect 64380 11364 64386 11416
rect 65320 11398 71858 11450
rect 71910 11398 71922 11450
rect 71974 11398 71986 11450
rect 72038 11398 72050 11450
rect 72102 11398 72114 11450
rect 72166 11398 74980 11450
rect 65320 11376 74980 11398
rect 63586 11296 63592 11348
rect 63644 11336 63650 11348
rect 63862 11336 63868 11348
rect 63644 11308 63868 11336
rect 63644 11296 63650 11308
rect 63862 11296 63868 11308
rect 63920 11296 63926 11348
rect 64966 11268 64972 11280
rect 63236 11240 64972 11268
rect 64966 11228 64972 11240
rect 65024 11228 65030 11280
rect 63402 11092 63408 11144
rect 63460 11132 63466 11144
rect 70854 11132 70860 11144
rect 63460 11104 70860 11132
rect 63460 11092 63466 11104
rect 70854 11092 70860 11104
rect 70912 11092 70918 11144
rect 65320 10906 74980 10928
rect 65320 10854 74210 10906
rect 74262 10854 74274 10906
rect 74326 10854 74338 10906
rect 74390 10854 74402 10906
rect 74454 10854 74466 10906
rect 74518 10854 74980 10906
rect 65320 10832 74980 10854
rect 63236 10452 63264 10570
rect 64874 10548 64880 10600
rect 64932 10588 64938 10600
rect 65610 10588 65616 10600
rect 64932 10560 65616 10588
rect 64932 10548 64938 10560
rect 65610 10548 65616 10560
rect 65668 10548 65674 10600
rect 65610 10452 65616 10464
rect 63236 10424 65616 10452
rect 65610 10412 65616 10424
rect 65668 10412 65674 10464
rect 65320 10362 74980 10384
rect 63494 10332 63500 10344
rect 63250 10304 63500 10332
rect 63494 10292 63500 10304
rect 63552 10292 63558 10344
rect 65320 10310 71858 10362
rect 71910 10310 71922 10362
rect 71974 10310 71986 10362
rect 72038 10310 72050 10362
rect 72102 10310 72114 10362
rect 72166 10310 74980 10362
rect 65320 10288 74980 10310
rect 65320 9818 74980 9840
rect 65320 9766 74210 9818
rect 74262 9766 74274 9818
rect 74326 9766 74338 9818
rect 74390 9766 74402 9818
rect 74454 9766 74466 9818
rect 74518 9766 74980 9818
rect 65320 9744 74980 9766
rect 64966 9364 64972 9376
rect 63236 9336 64972 9364
rect 64966 9324 64972 9336
rect 65024 9324 65030 9376
rect 65320 9274 74980 9296
rect 65320 9222 71858 9274
rect 71910 9222 71922 9274
rect 71974 9222 71986 9274
rect 72038 9222 72050 9274
rect 72102 9222 72114 9274
rect 72166 9222 74980 9274
rect 65320 9200 74980 9222
rect 65320 8730 74980 8752
rect 65320 8678 74210 8730
rect 74262 8678 74274 8730
rect 74326 8678 74338 8730
rect 74390 8678 74402 8730
rect 74454 8678 74466 8730
rect 74518 8678 74980 8730
rect 65320 8656 74980 8678
rect 65320 8186 74980 8208
rect 65320 8134 71858 8186
rect 71910 8134 71922 8186
rect 71974 8134 71986 8186
rect 72038 8134 72050 8186
rect 72102 8134 72114 8186
rect 72166 8134 74980 8186
rect 65320 8112 74980 8134
rect 67542 8072 67548 8084
rect 63144 8044 67548 8072
rect 59178 7828 59184 7880
rect 59236 7868 59242 7880
rect 63144 7868 63172 8044
rect 67542 8032 67548 8044
rect 67600 8032 67606 8084
rect 66806 8004 66812 8016
rect 63328 7976 66812 8004
rect 59236 7840 63172 7868
rect 59236 7828 59242 7840
rect 63218 7828 63224 7880
rect 63276 7868 63282 7880
rect 63328 7868 63356 7976
rect 66806 7964 66812 7976
rect 66864 7964 66870 8016
rect 63276 7840 63356 7868
rect 63276 7828 63282 7840
rect 64874 7828 64880 7880
rect 64932 7868 64938 7880
rect 65150 7868 65156 7880
rect 64932 7840 65156 7868
rect 64932 7828 64938 7840
rect 65150 7828 65156 7840
rect 65208 7828 65214 7880
rect 47302 7760 47308 7812
rect 47360 7800 47366 7812
rect 55766 7800 55772 7812
rect 47360 7772 55772 7800
rect 47360 7760 47366 7772
rect 55766 7760 55772 7772
rect 55824 7760 55830 7812
rect 59554 7760 59560 7812
rect 59612 7800 59618 7812
rect 63402 7800 63408 7812
rect 59612 7772 63408 7800
rect 59612 7760 59618 7772
rect 63402 7760 63408 7772
rect 63460 7760 63466 7812
rect 66346 7800 66352 7812
rect 63512 7772 66352 7800
rect 44818 7692 44824 7744
rect 44876 7732 44882 7744
rect 63512 7732 63540 7772
rect 66346 7760 66352 7772
rect 66404 7760 66410 7812
rect 44876 7704 63540 7732
rect 44876 7692 44882 7704
rect 65150 7692 65156 7744
rect 65208 7732 65214 7744
rect 65334 7732 65340 7744
rect 65208 7704 65340 7732
rect 65208 7692 65214 7704
rect 65334 7692 65340 7704
rect 65392 7692 65398 7744
rect 65320 7642 74980 7664
rect 33042 7556 33048 7608
rect 33100 7596 33106 7608
rect 63586 7596 63592 7608
rect 33100 7568 63592 7596
rect 33100 7556 33106 7568
rect 63586 7556 63592 7568
rect 63644 7556 63650 7608
rect 65320 7590 74210 7642
rect 74262 7590 74274 7642
rect 74326 7590 74338 7642
rect 74390 7590 74402 7642
rect 74454 7590 74466 7642
rect 74518 7590 74980 7642
rect 65320 7568 74980 7590
rect 67174 7528 67180 7540
rect 60706 7500 67180 7528
rect 55766 7420 55772 7472
rect 55824 7460 55830 7472
rect 60706 7460 60734 7500
rect 67174 7488 67180 7500
rect 67232 7488 67238 7540
rect 55824 7432 60734 7460
rect 55824 7420 55830 7432
rect 63126 7420 63132 7472
rect 63184 7460 63190 7472
rect 65794 7460 65800 7472
rect 63184 7432 65800 7460
rect 63184 7420 63190 7432
rect 65794 7420 65800 7432
rect 65852 7420 65858 7472
rect 62666 7352 62672 7404
rect 62724 7392 62730 7404
rect 67450 7392 67456 7404
rect 62724 7364 67456 7392
rect 62724 7352 62730 7364
rect 67450 7352 67456 7364
rect 67508 7352 67514 7404
rect 62298 7284 62304 7336
rect 62356 7324 62362 7336
rect 66070 7324 66076 7336
rect 62356 7296 66076 7324
rect 62356 7284 62362 7296
rect 66070 7284 66076 7296
rect 66128 7284 66134 7336
rect 55030 7216 55036 7268
rect 55088 7256 55094 7268
rect 64230 7256 64236 7268
rect 55088 7228 64236 7256
rect 55088 7216 55094 7228
rect 64230 7216 64236 7228
rect 64288 7216 64294 7268
rect 62758 7148 62764 7200
rect 62816 7188 62822 7200
rect 68738 7188 68744 7200
rect 62816 7160 68744 7188
rect 62816 7148 62822 7160
rect 68738 7148 68744 7160
rect 68796 7148 68802 7200
rect 65320 7098 74980 7120
rect 58618 7012 58624 7064
rect 58676 7052 58682 7064
rect 64506 7052 64512 7064
rect 58676 7024 64512 7052
rect 58676 7012 58682 7024
rect 64506 7012 64512 7024
rect 64564 7012 64570 7064
rect 65320 7046 71858 7098
rect 71910 7046 71922 7098
rect 71974 7046 71986 7098
rect 72038 7046 72050 7098
rect 72102 7046 72114 7098
rect 72166 7046 74980 7098
rect 65320 7024 74980 7046
rect 63310 6944 63316 6996
rect 63368 6984 63374 6996
rect 67910 6984 67916 6996
rect 63368 6956 67916 6984
rect 63368 6944 63374 6956
rect 67910 6944 67916 6956
rect 67968 6944 67974 6996
rect 61470 6876 61476 6928
rect 61528 6916 61534 6928
rect 63494 6916 63500 6928
rect 61528 6888 63500 6916
rect 61528 6876 61534 6888
rect 63494 6876 63500 6888
rect 63552 6876 63558 6928
rect 49050 6808 49056 6860
rect 49108 6848 49114 6860
rect 49108 6820 55904 6848
rect 49108 6808 49114 6820
rect 49786 6740 49792 6792
rect 49844 6780 49850 6792
rect 55766 6780 55772 6792
rect 49844 6752 55772 6780
rect 49844 6740 49850 6752
rect 55766 6740 55772 6752
rect 55824 6740 55830 6792
rect 55876 6780 55904 6820
rect 56502 6808 56508 6860
rect 56560 6848 56566 6860
rect 70394 6848 70400 6860
rect 56560 6820 70400 6848
rect 56560 6808 56566 6820
rect 70394 6808 70400 6820
rect 70452 6808 70458 6860
rect 66898 6780 66904 6792
rect 55876 6752 66904 6780
rect 66898 6740 66904 6752
rect 66956 6740 66962 6792
rect 66714 6712 66720 6724
rect 55876 6684 66720 6712
rect 47762 6604 47768 6656
rect 47820 6644 47826 6656
rect 55876 6644 55904 6684
rect 66714 6672 66720 6684
rect 66772 6672 66778 6724
rect 47820 6616 55904 6644
rect 47820 6604 47826 6616
rect 55950 6604 55956 6656
rect 56008 6644 56014 6656
rect 60918 6644 60924 6656
rect 56008 6616 60924 6644
rect 56008 6604 56014 6616
rect 60918 6604 60924 6616
rect 60976 6604 60982 6656
rect 61102 6604 61108 6656
rect 61160 6644 61166 6656
rect 68922 6644 68928 6656
rect 61160 6616 68928 6644
rect 61160 6604 61166 6616
rect 68922 6604 68928 6616
rect 68980 6604 68986 6656
rect 49602 6536 49608 6588
rect 49660 6576 49666 6588
rect 62758 6576 62764 6588
rect 49660 6548 62764 6576
rect 49660 6536 49666 6548
rect 62758 6536 62764 6548
rect 62816 6536 62822 6588
rect 65320 6554 74980 6576
rect 36722 6468 36728 6520
rect 36780 6508 36786 6520
rect 63126 6508 63132 6520
rect 36780 6480 63132 6508
rect 36780 6468 36786 6480
rect 63126 6468 63132 6480
rect 63184 6468 63190 6520
rect 65320 6502 74210 6554
rect 74262 6502 74274 6554
rect 74326 6502 74338 6554
rect 74390 6502 74402 6554
rect 74454 6502 74466 6554
rect 74518 6502 74980 6554
rect 65320 6480 74980 6502
rect 48222 6400 48228 6452
rect 48280 6440 48286 6452
rect 68002 6440 68008 6452
rect 48280 6412 64736 6440
rect 48280 6400 48286 6412
rect 46750 6332 46756 6384
rect 46808 6372 46814 6384
rect 61102 6372 61108 6384
rect 46808 6344 61108 6372
rect 46808 6332 46814 6344
rect 61102 6332 61108 6344
rect 61160 6332 61166 6384
rect 64708 6372 64736 6412
rect 64892 6412 68008 6440
rect 64892 6372 64920 6412
rect 68002 6400 68008 6412
rect 68060 6400 68066 6452
rect 63512 6344 64644 6372
rect 64708 6344 64920 6372
rect 42242 6264 42248 6316
rect 42300 6304 42306 6316
rect 63512 6304 63540 6344
rect 42300 6276 63540 6304
rect 64616 6304 64644 6344
rect 65794 6332 65800 6384
rect 65852 6372 65858 6384
rect 69842 6372 69848 6384
rect 65852 6344 69848 6372
rect 65852 6332 65858 6344
rect 69842 6332 69848 6344
rect 69900 6332 69906 6384
rect 67358 6304 67364 6316
rect 64616 6276 67364 6304
rect 42300 6264 42306 6276
rect 67358 6264 67364 6276
rect 67416 6264 67422 6316
rect 50706 6196 50712 6248
rect 50764 6236 50770 6248
rect 63310 6236 63316 6248
rect 50764 6208 63316 6236
rect 50764 6196 50770 6208
rect 63310 6196 63316 6208
rect 63368 6196 63374 6248
rect 63586 6196 63592 6248
rect 63644 6236 63650 6248
rect 64322 6236 64328 6248
rect 63644 6208 64328 6236
rect 63644 6196 63650 6208
rect 64322 6196 64328 6208
rect 64380 6196 64386 6248
rect 56318 6128 56324 6180
rect 56376 6168 56382 6180
rect 64966 6168 64972 6180
rect 56376 6140 64972 6168
rect 56376 6128 56382 6140
rect 64966 6128 64972 6140
rect 65024 6128 65030 6180
rect 56226 6060 56232 6112
rect 56284 6100 56290 6112
rect 69198 6100 69204 6112
rect 56284 6072 69204 6100
rect 56284 6060 56290 6072
rect 69198 6060 69204 6072
rect 69256 6060 69262 6112
rect 1012 6010 74980 6032
rect 1012 5958 71858 6010
rect 71910 5958 71922 6010
rect 71974 5958 71986 6010
rect 72038 5958 72050 6010
rect 72102 5958 72114 6010
rect 72166 5958 74980 6010
rect 1012 5936 74980 5958
rect 39482 5856 39488 5908
rect 39540 5856 39546 5908
rect 41690 5856 41696 5908
rect 41748 5856 41754 5908
rect 49602 5856 49608 5908
rect 49660 5856 49666 5908
rect 50706 5856 50712 5908
rect 50764 5856 50770 5908
rect 53653 5899 53711 5905
rect 53653 5865 53665 5899
rect 53699 5896 53711 5899
rect 53699 5868 61056 5896
rect 53699 5865 53711 5868
rect 53653 5859 53711 5865
rect 40402 5788 40408 5840
rect 40460 5788 40466 5840
rect 41598 5788 41604 5840
rect 41656 5828 41662 5840
rect 61028 5828 61056 5868
rect 61102 5856 61108 5908
rect 61160 5896 61166 5908
rect 72234 5896 72240 5908
rect 61160 5868 72240 5896
rect 61160 5856 61166 5868
rect 72234 5856 72240 5868
rect 72292 5856 72298 5908
rect 71498 5828 71504 5840
rect 41656 5800 45600 5828
rect 41656 5788 41662 5800
rect 29273 5763 29331 5769
rect 29273 5729 29285 5763
rect 29319 5760 29331 5763
rect 32306 5760 32312 5772
rect 29319 5732 32312 5760
rect 29319 5729 29331 5732
rect 29273 5723 29331 5729
rect 32306 5720 32312 5732
rect 32364 5720 32370 5772
rect 36357 5763 36415 5769
rect 36357 5729 36369 5763
rect 36403 5760 36415 5763
rect 44726 5760 44732 5772
rect 36403 5732 44732 5760
rect 36403 5729 36415 5732
rect 36357 5723 36415 5729
rect 44726 5720 44732 5732
rect 44784 5720 44790 5772
rect 28902 5652 28908 5704
rect 28960 5652 28966 5704
rect 29089 5695 29147 5701
rect 29089 5661 29101 5695
rect 29135 5692 29147 5695
rect 29546 5692 29552 5704
rect 29135 5664 29552 5692
rect 29135 5661 29147 5664
rect 29089 5655 29147 5661
rect 29546 5652 29552 5664
rect 29604 5652 29610 5704
rect 29917 5695 29975 5701
rect 29917 5661 29929 5695
rect 29963 5692 29975 5695
rect 30374 5692 30380 5704
rect 29963 5664 30380 5692
rect 29963 5661 29975 5664
rect 29917 5655 29975 5661
rect 30374 5652 30380 5664
rect 30432 5652 30438 5704
rect 30653 5695 30711 5701
rect 30653 5661 30665 5695
rect 30699 5692 30711 5695
rect 30742 5692 30748 5704
rect 30699 5664 30748 5692
rect 30699 5661 30711 5664
rect 30653 5655 30711 5661
rect 30742 5652 30748 5664
rect 30800 5652 30806 5704
rect 31386 5652 31392 5704
rect 31444 5652 31450 5704
rect 35158 5652 35164 5704
rect 35216 5692 35222 5704
rect 35713 5695 35771 5701
rect 35713 5692 35725 5695
rect 35216 5664 35725 5692
rect 35216 5652 35222 5664
rect 35713 5661 35725 5664
rect 35759 5661 35771 5695
rect 35713 5655 35771 5661
rect 36446 5652 36452 5704
rect 36504 5652 36510 5704
rect 36722 5652 36728 5704
rect 36780 5652 36786 5704
rect 37182 5652 37188 5704
rect 37240 5652 37246 5704
rect 38102 5652 38108 5704
rect 38160 5652 38166 5704
rect 38746 5652 38752 5704
rect 38804 5652 38810 5704
rect 38838 5652 38844 5704
rect 38896 5652 38902 5704
rect 39758 5652 39764 5704
rect 39816 5652 39822 5704
rect 40402 5652 40408 5704
rect 40460 5692 40466 5704
rect 41049 5695 41107 5701
rect 41049 5692 41061 5695
rect 40460 5664 41061 5692
rect 40460 5652 40466 5664
rect 41049 5661 41061 5664
rect 41095 5661 41107 5695
rect 41049 5655 41107 5661
rect 42702 5652 42708 5704
rect 42760 5652 42766 5704
rect 45572 5701 45600 5800
rect 51046 5800 60964 5828
rect 61028 5800 71504 5828
rect 46753 5763 46811 5769
rect 46753 5729 46765 5763
rect 46799 5760 46811 5763
rect 51046 5760 51074 5800
rect 46799 5732 51074 5760
rect 52181 5763 52239 5769
rect 46799 5729 46811 5732
rect 46753 5723 46811 5729
rect 52181 5729 52193 5763
rect 52227 5760 52239 5763
rect 60274 5760 60280 5772
rect 52227 5732 56456 5760
rect 52227 5729 52239 5732
rect 52181 5723 52239 5729
rect 45557 5695 45615 5701
rect 45557 5661 45569 5695
rect 45603 5661 45615 5695
rect 45557 5655 45615 5661
rect 47489 5695 47547 5701
rect 47489 5661 47501 5695
rect 47535 5661 47547 5695
rect 47489 5655 47547 5661
rect 29641 5627 29699 5633
rect 29641 5593 29653 5627
rect 29687 5624 29699 5627
rect 29687 5596 36676 5624
rect 29687 5593 29699 5596
rect 29641 5587 29699 5593
rect 29362 5516 29368 5568
rect 29420 5556 29426 5568
rect 30009 5559 30067 5565
rect 30009 5556 30021 5559
rect 29420 5528 30021 5556
rect 29420 5516 29426 5528
rect 30009 5525 30021 5528
rect 30055 5525 30067 5559
rect 30009 5519 30067 5525
rect 30834 5516 30840 5568
rect 30892 5516 30898 5568
rect 36648 5556 36676 5596
rect 38930 5584 38936 5636
rect 38988 5624 38994 5636
rect 47504 5624 47532 5655
rect 48958 5652 48964 5704
rect 49016 5652 49022 5704
rect 49694 5652 49700 5704
rect 49752 5692 49758 5704
rect 50065 5695 50123 5701
rect 50065 5692 50077 5695
rect 49752 5664 50077 5692
rect 49752 5652 49758 5664
rect 50065 5661 50077 5664
rect 50111 5661 50123 5695
rect 50065 5655 50123 5661
rect 50798 5652 50804 5704
rect 50856 5652 50862 5704
rect 51534 5652 51540 5704
rect 51592 5652 51598 5704
rect 52454 5652 52460 5704
rect 52512 5692 52518 5704
rect 53009 5695 53067 5701
rect 53009 5692 53021 5695
rect 52512 5664 53021 5692
rect 52512 5652 52518 5664
rect 53009 5661 53021 5664
rect 53055 5661 53067 5695
rect 53009 5655 53067 5661
rect 53834 5652 53840 5704
rect 53892 5692 53898 5704
rect 54389 5695 54447 5701
rect 54389 5692 54401 5695
rect 53892 5664 54401 5692
rect 53892 5652 53898 5664
rect 54389 5661 54401 5664
rect 54435 5661 54447 5695
rect 54389 5655 54447 5661
rect 55030 5652 55036 5704
rect 55088 5652 55094 5704
rect 55217 5695 55275 5701
rect 55217 5661 55229 5695
rect 55263 5661 55275 5695
rect 55217 5655 55275 5661
rect 38988 5596 47532 5624
rect 48685 5627 48743 5633
rect 38988 5584 38994 5596
rect 48685 5593 48697 5627
rect 48731 5624 48743 5627
rect 55232 5624 55260 5655
rect 56318 5652 56324 5704
rect 56376 5652 56382 5704
rect 56428 5692 56456 5732
rect 59832 5732 60280 5760
rect 56428 5664 56640 5692
rect 48731 5596 55260 5624
rect 56612 5624 56640 5664
rect 56686 5652 56692 5704
rect 56744 5652 56750 5704
rect 57333 5695 57391 5701
rect 57333 5661 57345 5695
rect 57379 5692 57391 5695
rect 59357 5695 59415 5701
rect 59357 5692 59369 5695
rect 57379 5664 59369 5692
rect 57379 5661 57391 5664
rect 57333 5655 57391 5661
rect 59357 5661 59369 5664
rect 59403 5661 59415 5695
rect 59357 5655 59415 5661
rect 59832 5624 59860 5732
rect 60274 5720 60280 5732
rect 60332 5720 60338 5772
rect 60458 5720 60464 5772
rect 60516 5720 60522 5772
rect 60936 5692 60964 5800
rect 71498 5788 71504 5800
rect 71556 5788 71562 5840
rect 61013 5763 61071 5769
rect 61013 5729 61025 5763
rect 61059 5760 61071 5763
rect 61286 5760 61292 5772
rect 61059 5732 61292 5760
rect 61059 5729 61071 5732
rect 61013 5723 61071 5729
rect 61286 5720 61292 5732
rect 61344 5720 61350 5772
rect 61378 5720 61384 5772
rect 61436 5760 61442 5772
rect 69750 5760 69756 5772
rect 61436 5732 69756 5760
rect 61436 5720 61442 5732
rect 69750 5720 69756 5732
rect 69808 5720 69814 5772
rect 67634 5692 67640 5704
rect 60936 5664 67640 5692
rect 67634 5652 67640 5664
rect 67692 5652 67698 5704
rect 56612 5596 59860 5624
rect 48731 5593 48743 5596
rect 48685 5587 48743 5593
rect 60274 5584 60280 5636
rect 60332 5624 60338 5636
rect 69474 5624 69480 5636
rect 60332 5596 69480 5624
rect 60332 5584 60338 5596
rect 69474 5584 69480 5596
rect 69532 5584 69538 5636
rect 37274 5556 37280 5568
rect 36648 5528 37280 5556
rect 37274 5516 37280 5528
rect 37332 5516 37338 5568
rect 37829 5559 37887 5565
rect 37829 5525 37841 5559
rect 37875 5556 37887 5559
rect 45462 5556 45468 5568
rect 37875 5528 45468 5556
rect 37875 5525 37887 5528
rect 37829 5519 37887 5525
rect 45462 5516 45468 5528
rect 45520 5516 45526 5568
rect 51445 5559 51503 5565
rect 51445 5525 51457 5559
rect 51491 5556 51503 5559
rect 58526 5556 58532 5568
rect 51491 5528 58532 5556
rect 51491 5525 51503 5528
rect 51445 5519 51503 5525
rect 58526 5516 58532 5528
rect 58584 5516 58590 5568
rect 60001 5559 60059 5565
rect 60001 5525 60013 5559
rect 60047 5556 60059 5559
rect 66162 5556 66168 5568
rect 60047 5528 66168 5556
rect 60047 5525 60059 5528
rect 60001 5519 60059 5525
rect 66162 5516 66168 5528
rect 66220 5516 66226 5568
rect 69934 5516 69940 5568
rect 69992 5556 69998 5568
rect 71130 5556 71136 5568
rect 69992 5528 71136 5556
rect 69992 5516 69998 5528
rect 71130 5516 71136 5528
rect 71188 5516 71194 5568
rect 71590 5516 71596 5568
rect 71648 5556 71654 5568
rect 73430 5556 73436 5568
rect 71648 5528 73436 5556
rect 71648 5516 71654 5528
rect 73430 5516 73436 5528
rect 73488 5516 73494 5568
rect 1012 5466 74980 5488
rect 1012 5414 4210 5466
rect 4262 5414 4274 5466
rect 4326 5414 4338 5466
rect 4390 5414 4402 5466
rect 4454 5414 4466 5466
rect 4518 5414 14210 5466
rect 14262 5414 14274 5466
rect 14326 5414 14338 5466
rect 14390 5414 14402 5466
rect 14454 5414 14466 5466
rect 14518 5414 24210 5466
rect 24262 5414 24274 5466
rect 24326 5414 24338 5466
rect 24390 5414 24402 5466
rect 24454 5414 24466 5466
rect 24518 5414 34210 5466
rect 34262 5414 34274 5466
rect 34326 5414 34338 5466
rect 34390 5414 34402 5466
rect 34454 5414 34466 5466
rect 34518 5414 44210 5466
rect 44262 5414 44274 5466
rect 44326 5414 44338 5466
rect 44390 5414 44402 5466
rect 44454 5414 44466 5466
rect 44518 5414 54210 5466
rect 54262 5414 54274 5466
rect 54326 5414 54338 5466
rect 54390 5414 54402 5466
rect 54454 5414 54466 5466
rect 54518 5414 64210 5466
rect 64262 5414 64274 5466
rect 64326 5414 64338 5466
rect 64390 5414 64402 5466
rect 64454 5414 64466 5466
rect 64518 5414 74210 5466
rect 74262 5414 74274 5466
rect 74326 5414 74338 5466
rect 74390 5414 74402 5466
rect 74454 5414 74466 5466
rect 74518 5414 74980 5466
rect 1012 5392 74980 5414
rect 35713 5355 35771 5361
rect 35713 5321 35725 5355
rect 35759 5352 35771 5355
rect 36446 5352 36452 5364
rect 35759 5324 36452 5352
rect 35759 5321 35771 5324
rect 35713 5315 35771 5321
rect 36446 5312 36452 5324
rect 36504 5312 36510 5364
rect 37829 5355 37887 5361
rect 37829 5321 37841 5355
rect 37875 5352 37887 5355
rect 41598 5352 41604 5364
rect 37875 5324 41604 5352
rect 37875 5321 37887 5324
rect 37829 5315 37887 5321
rect 41598 5312 41604 5324
rect 41656 5312 41662 5364
rect 42153 5355 42211 5361
rect 42153 5321 42165 5355
rect 42199 5352 42211 5355
rect 42199 5324 42288 5352
rect 42199 5321 42211 5324
rect 42153 5315 42211 5321
rect 42260 5296 42288 5324
rect 42702 5312 42708 5364
rect 42760 5352 42766 5364
rect 42797 5355 42855 5361
rect 42797 5352 42809 5355
rect 42760 5324 42809 5352
rect 42760 5312 42766 5324
rect 42797 5321 42809 5324
rect 42843 5321 42855 5355
rect 42797 5315 42855 5321
rect 42886 5312 42892 5364
rect 42944 5352 42950 5364
rect 42944 5324 46244 5352
rect 42944 5312 42950 5324
rect 28905 5287 28963 5293
rect 28905 5253 28917 5287
rect 28951 5284 28963 5287
rect 38102 5284 38108 5296
rect 28951 5256 38108 5284
rect 28951 5253 28963 5256
rect 28905 5247 28963 5253
rect 38102 5244 38108 5256
rect 38160 5244 38166 5296
rect 42242 5244 42248 5296
rect 42300 5244 42306 5296
rect 46106 5244 46112 5296
rect 46164 5244 46170 5296
rect 46216 5284 46244 5324
rect 47302 5312 47308 5364
rect 47360 5312 47366 5364
rect 48222 5312 48228 5364
rect 48280 5312 48286 5364
rect 49050 5312 49056 5364
rect 49108 5312 49114 5364
rect 49786 5312 49792 5364
rect 49844 5312 49850 5364
rect 50525 5355 50583 5361
rect 50525 5321 50537 5355
rect 50571 5352 50583 5355
rect 53466 5352 53472 5364
rect 50571 5324 53472 5352
rect 50571 5321 50583 5324
rect 50525 5315 50583 5321
rect 53466 5312 53472 5324
rect 53524 5312 53530 5364
rect 54018 5312 54024 5364
rect 54076 5312 54082 5364
rect 54757 5355 54815 5361
rect 54757 5321 54769 5355
rect 54803 5352 54815 5355
rect 56965 5355 57023 5361
rect 54803 5324 56916 5352
rect 54803 5321 54815 5324
rect 54757 5315 54815 5321
rect 48958 5284 48964 5296
rect 46216 5256 48964 5284
rect 48958 5244 48964 5256
rect 49016 5244 49022 5296
rect 51997 5287 52055 5293
rect 51997 5253 52009 5287
rect 52043 5284 52055 5287
rect 52043 5256 55720 5284
rect 52043 5253 52055 5256
rect 51997 5247 52055 5253
rect 29178 5176 29184 5228
rect 29236 5176 29242 5228
rect 29362 5176 29368 5228
rect 29420 5176 29426 5228
rect 32125 5219 32183 5225
rect 32125 5185 32137 5219
rect 32171 5216 32183 5219
rect 32214 5216 32220 5228
rect 32171 5188 32220 5216
rect 32171 5185 32183 5188
rect 32125 5179 32183 5185
rect 32214 5176 32220 5188
rect 32272 5176 32278 5228
rect 37274 5176 37280 5228
rect 37332 5216 37338 5228
rect 38565 5219 38623 5225
rect 38565 5216 38577 5219
rect 37332 5188 38577 5216
rect 37332 5176 37338 5188
rect 38565 5185 38577 5188
rect 38611 5185 38623 5219
rect 41509 5219 41567 5225
rect 41509 5216 41521 5219
rect 38565 5179 38623 5185
rect 38672 5188 41521 5216
rect 25038 5108 25044 5160
rect 25096 5148 25102 5160
rect 26053 5151 26111 5157
rect 26053 5148 26065 5151
rect 25096 5120 26065 5148
rect 25096 5108 25102 5120
rect 26053 5117 26065 5120
rect 26099 5117 26111 5151
rect 26053 5111 26111 5117
rect 26142 5108 26148 5160
rect 26200 5148 26206 5160
rect 27433 5151 27491 5157
rect 27433 5148 27445 5151
rect 26200 5120 27445 5148
rect 26200 5108 26206 5120
rect 27433 5117 27445 5120
rect 27479 5117 27491 5151
rect 27433 5111 27491 5117
rect 28350 5108 28356 5160
rect 28408 5148 28414 5160
rect 28445 5151 28503 5157
rect 28445 5148 28457 5151
rect 28408 5120 28457 5148
rect 28408 5108 28414 5120
rect 28445 5117 28457 5120
rect 28491 5117 28503 5151
rect 28445 5111 28503 5117
rect 29917 5151 29975 5157
rect 29917 5117 29929 5151
rect 29963 5148 29975 5151
rect 30009 5151 30067 5157
rect 30009 5148 30021 5151
rect 29963 5120 30021 5148
rect 29963 5117 29975 5120
rect 29917 5111 29975 5117
rect 30009 5117 30021 5120
rect 30055 5117 30067 5151
rect 30009 5111 30067 5117
rect 31113 5151 31171 5157
rect 31113 5117 31125 5151
rect 31159 5148 31171 5151
rect 31294 5148 31300 5160
rect 31159 5120 31300 5148
rect 31159 5117 31171 5120
rect 31113 5111 31171 5117
rect 31294 5108 31300 5120
rect 31352 5108 31358 5160
rect 33410 5108 33416 5160
rect 33468 5108 33474 5160
rect 33778 5108 33784 5160
rect 33836 5148 33842 5160
rect 35069 5151 35127 5157
rect 35069 5148 35081 5151
rect 33836 5120 35081 5148
rect 33836 5108 33842 5120
rect 35069 5117 35081 5120
rect 35115 5117 35127 5151
rect 35069 5111 35127 5117
rect 36538 5108 36544 5160
rect 36596 5148 36602 5160
rect 37185 5151 37243 5157
rect 37185 5148 37197 5151
rect 36596 5120 37197 5148
rect 36596 5108 36602 5120
rect 37185 5117 37197 5120
rect 37231 5117 37243 5151
rect 37185 5111 37243 5117
rect 37734 5108 37740 5160
rect 37792 5148 37798 5160
rect 38672 5148 38700 5188
rect 41509 5185 41521 5188
rect 41555 5185 41567 5219
rect 41509 5179 41567 5185
rect 44082 5176 44088 5228
rect 44140 5176 44146 5228
rect 44726 5176 44732 5228
rect 44784 5176 44790 5228
rect 45462 5176 45468 5228
rect 45520 5176 45526 5228
rect 46198 5176 46204 5228
rect 46256 5216 46262 5228
rect 52822 5216 52828 5228
rect 46256 5188 52828 5216
rect 46256 5176 46262 5188
rect 52822 5176 52828 5188
rect 52880 5176 52886 5228
rect 55692 5225 55720 5256
rect 55858 5244 55864 5296
rect 55916 5284 55922 5296
rect 56888 5284 56916 5324
rect 56965 5321 56977 5355
rect 57011 5352 57023 5355
rect 60366 5352 60372 5364
rect 57011 5324 60372 5352
rect 57011 5321 57023 5324
rect 56965 5315 57023 5321
rect 60366 5312 60372 5324
rect 60424 5312 60430 5364
rect 67726 5352 67732 5364
rect 60476 5324 67732 5352
rect 60476 5284 60504 5324
rect 67726 5312 67732 5324
rect 67784 5312 67790 5364
rect 55916 5256 56456 5284
rect 56888 5256 60504 5284
rect 55916 5244 55922 5256
rect 56428 5225 56456 5256
rect 60550 5244 60556 5296
rect 60608 5284 60614 5296
rect 69290 5284 69296 5296
rect 60608 5256 69296 5284
rect 60608 5244 60614 5256
rect 69290 5244 69296 5256
rect 69348 5244 69354 5296
rect 55677 5219 55735 5225
rect 55677 5185 55689 5219
rect 55723 5185 55735 5219
rect 55677 5179 55735 5185
rect 56413 5219 56471 5225
rect 56413 5185 56425 5219
rect 56459 5185 56471 5219
rect 56413 5179 56471 5185
rect 56594 5176 56600 5228
rect 56652 5216 56658 5228
rect 69106 5216 69112 5228
rect 56652 5188 69112 5216
rect 56652 5176 56658 5188
rect 69106 5176 69112 5188
rect 69164 5176 69170 5228
rect 37792 5120 38700 5148
rect 37792 5108 37798 5120
rect 39206 5108 39212 5160
rect 39264 5108 39270 5160
rect 40126 5108 40132 5160
rect 40184 5108 40190 5160
rect 46658 5108 46664 5160
rect 46716 5108 46722 5160
rect 47578 5108 47584 5160
rect 47636 5108 47642 5160
rect 48406 5108 48412 5160
rect 48464 5108 48470 5160
rect 49142 5108 49148 5160
rect 49200 5108 49206 5160
rect 49786 5108 49792 5160
rect 49844 5148 49850 5160
rect 49881 5151 49939 5157
rect 49881 5148 49893 5151
rect 49844 5120 49893 5148
rect 49844 5108 49850 5120
rect 49881 5117 49893 5120
rect 49927 5117 49939 5151
rect 49881 5111 49939 5117
rect 50154 5108 50160 5160
rect 50212 5148 50218 5160
rect 50617 5151 50675 5157
rect 50617 5148 50629 5151
rect 50212 5120 50629 5148
rect 50212 5108 50218 5120
rect 50617 5117 50629 5120
rect 50663 5117 50675 5151
rect 50617 5111 50675 5117
rect 51258 5108 51264 5160
rect 51316 5108 51322 5160
rect 51350 5108 51356 5160
rect 51408 5108 51414 5160
rect 51718 5108 51724 5160
rect 51776 5148 51782 5160
rect 52641 5151 52699 5157
rect 52641 5148 52653 5151
rect 51776 5120 52653 5148
rect 51776 5108 51782 5120
rect 52641 5117 52653 5120
rect 52687 5117 52699 5151
rect 52641 5111 52699 5117
rect 53282 5108 53288 5160
rect 53340 5108 53346 5160
rect 53374 5108 53380 5160
rect 53432 5108 53438 5160
rect 53466 5108 53472 5160
rect 53524 5148 53530 5160
rect 54113 5151 54171 5157
rect 54113 5148 54125 5151
rect 53524 5120 54125 5148
rect 53524 5108 53530 5120
rect 54113 5117 54125 5120
rect 54159 5117 54171 5151
rect 54113 5111 54171 5117
rect 54846 5108 54852 5160
rect 54904 5108 54910 5160
rect 55398 5108 55404 5160
rect 55456 5148 55462 5160
rect 69566 5148 69572 5160
rect 55456 5120 69572 5148
rect 55456 5108 55462 5120
rect 69566 5108 69572 5120
rect 69624 5108 69630 5160
rect 23566 5040 23572 5092
rect 23624 5080 23630 5092
rect 26881 5083 26939 5089
rect 26881 5080 26893 5083
rect 23624 5052 26893 5080
rect 23624 5040 23630 5052
rect 26881 5049 26893 5052
rect 26927 5049 26939 5083
rect 26881 5043 26939 5049
rect 32401 5083 32459 5089
rect 32401 5049 32413 5083
rect 32447 5080 32459 5083
rect 39942 5080 39948 5092
rect 32447 5052 39948 5080
rect 32447 5049 32459 5052
rect 32401 5043 32459 5049
rect 39942 5040 39948 5052
rect 40000 5040 40006 5092
rect 40773 5083 40831 5089
rect 40773 5049 40785 5083
rect 40819 5080 40831 5083
rect 43622 5080 43628 5092
rect 40819 5052 43628 5080
rect 40819 5049 40831 5052
rect 40773 5043 40831 5049
rect 43622 5040 43628 5052
rect 43680 5040 43686 5092
rect 69382 5080 69388 5092
rect 47228 5052 69388 5080
rect 26694 4972 26700 5024
rect 26752 4972 26758 5024
rect 27890 4972 27896 5024
rect 27948 4972 27954 5024
rect 30650 4972 30656 5024
rect 30708 4972 30714 5024
rect 31570 4972 31576 5024
rect 31628 5012 31634 5024
rect 31665 5015 31723 5021
rect 31665 5012 31677 5015
rect 31628 4984 31677 5012
rect 31628 4972 31634 4984
rect 31665 4981 31677 4984
rect 31711 4981 31723 5015
rect 31665 4975 31723 4981
rect 32858 4972 32864 5024
rect 32916 4972 32922 5024
rect 36078 4972 36084 5024
rect 36136 5012 36142 5024
rect 38838 5012 38844 5024
rect 36136 4984 38844 5012
rect 36136 4972 36142 4984
rect 38838 4972 38844 4984
rect 38896 4972 38902 5024
rect 45373 5015 45431 5021
rect 45373 4981 45385 5015
rect 45419 5012 45431 5015
rect 47228 5012 47256 5052
rect 69382 5040 69388 5052
rect 69440 5040 69446 5092
rect 45419 4984 47256 5012
rect 45419 4981 45431 4984
rect 45373 4975 45431 4981
rect 55490 4972 55496 5024
rect 55548 4972 55554 5024
rect 56226 4972 56232 5024
rect 56284 4972 56290 5024
rect 56410 4972 56416 5024
rect 56468 5012 56474 5024
rect 63218 5012 63224 5024
rect 56468 4984 63224 5012
rect 56468 4972 56474 4984
rect 63218 4972 63224 4984
rect 63276 4972 63282 5024
rect 1012 4922 74980 4944
rect 1012 4870 1858 4922
rect 1910 4870 1922 4922
rect 1974 4870 1986 4922
rect 2038 4870 2050 4922
rect 2102 4870 2114 4922
rect 2166 4870 11858 4922
rect 11910 4870 11922 4922
rect 11974 4870 11986 4922
rect 12038 4870 12050 4922
rect 12102 4870 12114 4922
rect 12166 4870 21858 4922
rect 21910 4870 21922 4922
rect 21974 4870 21986 4922
rect 22038 4870 22050 4922
rect 22102 4870 22114 4922
rect 22166 4870 31858 4922
rect 31910 4870 31922 4922
rect 31974 4870 31986 4922
rect 32038 4870 32050 4922
rect 32102 4870 32114 4922
rect 32166 4870 41858 4922
rect 41910 4870 41922 4922
rect 41974 4870 41986 4922
rect 42038 4870 42050 4922
rect 42102 4870 42114 4922
rect 42166 4870 51858 4922
rect 51910 4870 51922 4922
rect 51974 4870 51986 4922
rect 52038 4870 52050 4922
rect 52102 4870 52114 4922
rect 52166 4870 61858 4922
rect 61910 4870 61922 4922
rect 61974 4870 61986 4922
rect 62038 4870 62050 4922
rect 62102 4870 62114 4922
rect 62166 4870 71858 4922
rect 71910 4870 71922 4922
rect 71974 4870 71986 4922
rect 72038 4870 72050 4922
rect 72102 4870 72114 4922
rect 72166 4870 74980 4922
rect 1012 4848 74980 4870
rect 26142 4768 26148 4820
rect 26200 4768 26206 4820
rect 31294 4768 31300 4820
rect 31352 4768 31358 4820
rect 33778 4768 33784 4820
rect 33836 4768 33842 4820
rect 35529 4811 35587 4817
rect 35529 4777 35541 4811
rect 35575 4808 35587 4811
rect 42889 4811 42947 4817
rect 35575 4780 42288 4808
rect 35575 4777 35587 4780
rect 35529 4771 35587 4777
rect 26881 4743 26939 4749
rect 26881 4709 26893 4743
rect 26927 4740 26939 4743
rect 29546 4740 29552 4752
rect 26927 4712 29552 4740
rect 26927 4709 26939 4712
rect 26881 4703 26939 4709
rect 29546 4700 29552 4712
rect 29604 4700 29610 4752
rect 34440 4712 40540 4740
rect 25593 4675 25651 4681
rect 25593 4641 25605 4675
rect 25639 4672 25651 4675
rect 26326 4672 26332 4684
rect 25639 4644 26332 4672
rect 25639 4641 25651 4644
rect 25593 4635 25651 4641
rect 26326 4632 26332 4644
rect 26384 4632 26390 4684
rect 34440 4681 34468 4712
rect 28353 4675 28411 4681
rect 28353 4641 28365 4675
rect 28399 4672 28411 4675
rect 34425 4675 34483 4681
rect 28399 4644 34100 4672
rect 28399 4641 28411 4644
rect 28353 4635 28411 4641
rect 24854 4564 24860 4616
rect 24912 4604 24918 4616
rect 25041 4607 25099 4613
rect 25041 4604 25053 4607
rect 24912 4576 25053 4604
rect 24912 4564 24918 4576
rect 25041 4573 25053 4576
rect 25087 4573 25099 4607
rect 25041 4567 25099 4573
rect 26234 4564 26240 4616
rect 26292 4564 26298 4616
rect 27985 4607 28043 4613
rect 27985 4573 27997 4607
rect 28031 4604 28043 4607
rect 28074 4604 28080 4616
rect 28031 4576 28080 4604
rect 28031 4573 28043 4576
rect 27985 4567 28043 4573
rect 28074 4564 28080 4576
rect 28132 4564 28138 4616
rect 28537 4607 28595 4613
rect 28537 4573 28549 4607
rect 28583 4573 28595 4607
rect 28537 4567 28595 4573
rect 28552 4536 28580 4567
rect 28626 4564 28632 4616
rect 28684 4564 28690 4616
rect 29822 4564 29828 4616
rect 29880 4564 29886 4616
rect 31205 4607 31263 4613
rect 31205 4573 31217 4607
rect 31251 4604 31263 4607
rect 31294 4604 31300 4616
rect 31251 4576 31300 4604
rect 31251 4573 31263 4576
rect 31205 4567 31263 4573
rect 31294 4564 31300 4576
rect 31352 4564 31358 4616
rect 31849 4607 31907 4613
rect 31849 4573 31861 4607
rect 31895 4573 31907 4607
rect 31849 4567 31907 4573
rect 29638 4536 29644 4548
rect 28552 4508 29644 4536
rect 29638 4496 29644 4508
rect 29696 4496 29702 4548
rect 30926 4496 30932 4548
rect 30984 4536 30990 4548
rect 31864 4536 31892 4567
rect 32674 4564 32680 4616
rect 32732 4604 32738 4616
rect 32953 4607 33011 4613
rect 32953 4604 32965 4607
rect 32732 4576 32965 4604
rect 32732 4564 32738 4576
rect 32953 4573 32965 4576
rect 32999 4573 33011 4607
rect 32953 4567 33011 4573
rect 33134 4564 33140 4616
rect 33192 4564 33198 4616
rect 33962 4564 33968 4616
rect 34020 4564 34026 4616
rect 34072 4604 34100 4644
rect 34425 4641 34437 4675
rect 34471 4641 34483 4675
rect 36078 4672 36084 4684
rect 34425 4635 34483 4641
rect 34532 4644 36084 4672
rect 34532 4604 34560 4644
rect 36078 4632 36084 4644
rect 36136 4632 36142 4684
rect 36173 4675 36231 4681
rect 36173 4641 36185 4675
rect 36219 4672 36231 4675
rect 40512 4672 40540 4712
rect 40586 4700 40592 4752
rect 40644 4700 40650 4752
rect 40696 4712 42196 4740
rect 40696 4672 40724 4712
rect 36219 4644 37872 4672
rect 40512 4644 40724 4672
rect 36219 4641 36231 4644
rect 36173 4635 36231 4641
rect 34072 4576 34560 4604
rect 34606 4564 34612 4616
rect 34664 4564 34670 4616
rect 34885 4607 34943 4613
rect 34885 4573 34897 4607
rect 34931 4604 34943 4607
rect 34931 4576 35894 4604
rect 34931 4573 34943 4576
rect 34885 4567 34943 4573
rect 30984 4508 31892 4536
rect 30984 4496 30990 4508
rect 35250 4496 35256 4548
rect 35308 4496 35314 4548
rect 35866 4536 35894 4576
rect 36354 4564 36360 4616
rect 36412 4564 36418 4616
rect 37734 4604 37740 4616
rect 36464 4576 37740 4604
rect 36464 4536 36492 4576
rect 37734 4564 37740 4576
rect 37792 4564 37798 4616
rect 37844 4604 37872 4644
rect 37844 4576 39528 4604
rect 35866 4508 36492 4536
rect 36817 4539 36875 4545
rect 36817 4505 36829 4539
rect 36863 4536 36875 4539
rect 36906 4536 36912 4548
rect 36863 4508 36912 4536
rect 36863 4505 36875 4508
rect 36817 4499 36875 4505
rect 36906 4496 36912 4508
rect 36964 4496 36970 4548
rect 38010 4496 38016 4548
rect 38068 4496 38074 4548
rect 39500 4536 39528 4576
rect 39942 4564 39948 4616
rect 40000 4564 40006 4616
rect 40218 4564 40224 4616
rect 40276 4604 40282 4616
rect 41325 4607 41383 4613
rect 41325 4604 41337 4607
rect 40276 4576 41337 4604
rect 40276 4564 40282 4576
rect 41325 4573 41337 4576
rect 41371 4573 41383 4607
rect 42168 4604 42196 4712
rect 42260 4681 42288 4780
rect 42889 4777 42901 4811
rect 42935 4808 42947 4811
rect 49142 4808 49148 4820
rect 42935 4780 49148 4808
rect 42935 4777 42947 4780
rect 42889 4771 42947 4777
rect 49142 4768 49148 4780
rect 49200 4768 49206 4820
rect 54018 4768 54024 4820
rect 54076 4808 54082 4820
rect 65702 4808 65708 4820
rect 54076 4780 65708 4808
rect 54076 4768 54082 4780
rect 65702 4768 65708 4780
rect 65760 4768 65766 4820
rect 43622 4700 43628 4752
rect 43680 4740 43686 4752
rect 66438 4740 66444 4752
rect 43680 4712 66444 4740
rect 43680 4700 43686 4712
rect 66438 4700 66444 4712
rect 66496 4700 66502 4752
rect 42245 4675 42303 4681
rect 42245 4641 42257 4675
rect 42291 4641 42303 4675
rect 67266 4672 67272 4684
rect 42245 4635 42303 4641
rect 42352 4644 67272 4672
rect 42352 4604 42380 4644
rect 67266 4632 67272 4644
rect 67324 4632 67330 4684
rect 42168 4576 42380 4604
rect 42981 4607 43039 4613
rect 41325 4567 41383 4573
rect 42981 4573 42993 4607
rect 43027 4573 43039 4607
rect 42981 4567 43039 4573
rect 42996 4536 43024 4567
rect 44082 4564 44088 4616
rect 44140 4564 44146 4616
rect 44729 4607 44787 4613
rect 44729 4573 44741 4607
rect 44775 4604 44787 4607
rect 44818 4604 44824 4616
rect 44775 4576 44824 4604
rect 44775 4573 44787 4576
rect 44729 4567 44787 4573
rect 44818 4564 44824 4576
rect 44876 4564 44882 4616
rect 45002 4564 45008 4616
rect 45060 4564 45066 4616
rect 45094 4564 45100 4616
rect 45152 4604 45158 4616
rect 46109 4607 46167 4613
rect 46109 4604 46121 4607
rect 45152 4576 46121 4604
rect 45152 4564 45158 4576
rect 46109 4573 46121 4576
rect 46155 4573 46167 4607
rect 46109 4567 46167 4573
rect 46750 4564 46756 4616
rect 46808 4564 46814 4616
rect 47210 4564 47216 4616
rect 47268 4564 47274 4616
rect 47762 4564 47768 4616
rect 47820 4564 47826 4616
rect 47854 4564 47860 4616
rect 47912 4564 47918 4616
rect 49602 4564 49608 4616
rect 49660 4604 49666 4616
rect 51169 4607 51227 4613
rect 51169 4604 51181 4607
rect 49660 4576 51181 4604
rect 49660 4564 49666 4576
rect 51169 4573 51181 4576
rect 51215 4573 51227 4607
rect 51169 4567 51227 4573
rect 53282 4564 53288 4616
rect 53340 4604 53346 4616
rect 60550 4604 60556 4616
rect 53340 4576 60556 4604
rect 53340 4564 53346 4576
rect 60550 4564 60556 4576
rect 60608 4564 60614 4616
rect 39500 4508 43024 4536
rect 43625 4539 43683 4545
rect 43625 4505 43637 4539
rect 43671 4536 43683 4539
rect 66530 4536 66536 4548
rect 43671 4508 66536 4536
rect 43671 4505 43683 4508
rect 43625 4499 43683 4505
rect 66530 4496 66536 4508
rect 66588 4496 66594 4548
rect 23474 4428 23480 4480
rect 23532 4468 23538 4480
rect 24489 4471 24547 4477
rect 24489 4468 24501 4471
rect 23532 4440 24501 4468
rect 23532 4428 23538 4440
rect 24489 4437 24501 4440
rect 24535 4437 24547 4471
rect 24489 4431 24547 4437
rect 27338 4428 27344 4480
rect 27396 4428 27402 4480
rect 29270 4428 29276 4480
rect 29328 4428 29334 4480
rect 30466 4428 30472 4480
rect 30524 4428 30530 4480
rect 30558 4428 30564 4480
rect 30616 4428 30622 4480
rect 32398 4428 32404 4480
rect 32456 4428 32462 4480
rect 36722 4428 36728 4480
rect 36780 4428 36786 4480
rect 37918 4428 37924 4480
rect 37976 4428 37982 4480
rect 41969 4471 42027 4477
rect 41969 4437 41981 4471
rect 42015 4468 42027 4471
rect 42886 4468 42892 4480
rect 42015 4440 42892 4468
rect 42015 4437 42027 4440
rect 41969 4431 42027 4437
rect 42886 4428 42892 4440
rect 42944 4428 42950 4480
rect 45646 4428 45652 4480
rect 45704 4428 45710 4480
rect 48501 4471 48559 4477
rect 48501 4437 48513 4471
rect 48547 4468 48559 4471
rect 51718 4468 51724 4480
rect 48547 4440 51724 4468
rect 48547 4437 48559 4440
rect 48501 4431 48559 4437
rect 51718 4428 51724 4440
rect 51776 4428 51782 4480
rect 51813 4471 51871 4477
rect 51813 4437 51825 4471
rect 51859 4468 51871 4471
rect 56686 4468 56692 4480
rect 51859 4440 56692 4468
rect 51859 4437 51871 4440
rect 51813 4431 51871 4437
rect 56686 4428 56692 4440
rect 56744 4428 56750 4480
rect 1012 4378 74980 4400
rect 1012 4326 4210 4378
rect 4262 4326 4274 4378
rect 4326 4326 4338 4378
rect 4390 4326 4402 4378
rect 4454 4326 4466 4378
rect 4518 4326 14210 4378
rect 14262 4326 14274 4378
rect 14326 4326 14338 4378
rect 14390 4326 14402 4378
rect 14454 4326 14466 4378
rect 14518 4326 24210 4378
rect 24262 4326 24274 4378
rect 24326 4326 24338 4378
rect 24390 4326 24402 4378
rect 24454 4326 24466 4378
rect 24518 4326 34210 4378
rect 34262 4326 34274 4378
rect 34326 4326 34338 4378
rect 34390 4326 34402 4378
rect 34454 4326 34466 4378
rect 34518 4326 44210 4378
rect 44262 4326 44274 4378
rect 44326 4326 44338 4378
rect 44390 4326 44402 4378
rect 44454 4326 44466 4378
rect 44518 4326 54210 4378
rect 54262 4326 54274 4378
rect 54326 4326 54338 4378
rect 54390 4326 54402 4378
rect 54454 4326 54466 4378
rect 54518 4326 64210 4378
rect 64262 4326 64274 4378
rect 64326 4326 64338 4378
rect 64390 4326 64402 4378
rect 64454 4326 64466 4378
rect 64518 4326 74210 4378
rect 74262 4326 74274 4378
rect 74326 4326 74338 4378
rect 74390 4326 74402 4378
rect 74454 4326 74466 4378
rect 74518 4326 74980 4378
rect 1012 4304 74980 4326
rect 36722 4224 36728 4276
rect 36780 4264 36786 4276
rect 43530 4264 43536 4276
rect 36780 4236 43536 4264
rect 36780 4224 36786 4236
rect 43530 4224 43536 4236
rect 43588 4224 43594 4276
rect 45646 4224 45652 4276
rect 45704 4264 45710 4276
rect 56410 4264 56416 4276
rect 45704 4236 56416 4264
rect 45704 4224 45710 4236
rect 56410 4224 56416 4236
rect 56468 4224 56474 4276
rect 60458 4224 60464 4276
rect 60516 4264 60522 4276
rect 63862 4264 63868 4276
rect 60516 4236 63868 4264
rect 60516 4224 60522 4236
rect 63862 4224 63868 4236
rect 63920 4224 63926 4276
rect 31110 4156 31116 4208
rect 31168 4196 31174 4208
rect 32858 4196 32864 4208
rect 31168 4168 32864 4196
rect 31168 4156 31174 4168
rect 32858 4156 32864 4168
rect 32916 4156 32922 4208
rect 37918 4156 37924 4208
rect 37976 4196 37982 4208
rect 37976 4168 44312 4196
rect 37976 4156 37982 4168
rect 26510 4088 26516 4140
rect 26568 4128 26574 4140
rect 26881 4131 26939 4137
rect 26881 4128 26893 4131
rect 26568 4100 26893 4128
rect 26568 4088 26574 4100
rect 26881 4097 26893 4100
rect 26927 4097 26939 4131
rect 26881 4091 26939 4097
rect 27525 4131 27583 4137
rect 27525 4097 27537 4131
rect 27571 4128 27583 4131
rect 28905 4131 28963 4137
rect 27571 4100 28856 4128
rect 27571 4097 27583 4100
rect 27525 4091 27583 4097
rect 24578 4020 24584 4072
rect 24636 4020 24642 4072
rect 25130 4020 25136 4072
rect 25188 4060 25194 4072
rect 25869 4063 25927 4069
rect 25869 4060 25881 4063
rect 25188 4032 25881 4060
rect 25188 4020 25194 4032
rect 25869 4029 25881 4032
rect 25915 4029 25927 4063
rect 25869 4023 25927 4029
rect 25958 4020 25964 4072
rect 26016 4060 26022 4072
rect 26605 4063 26663 4069
rect 26605 4060 26617 4063
rect 26016 4032 26617 4060
rect 26016 4020 26022 4032
rect 26605 4029 26617 4032
rect 26651 4029 26663 4063
rect 26605 4023 26663 4029
rect 27157 4063 27215 4069
rect 27157 4029 27169 4063
rect 27203 4029 27215 4063
rect 27157 4023 27215 4029
rect 27172 3992 27200 4023
rect 27706 4020 27712 4072
rect 27764 4060 27770 4072
rect 28169 4063 28227 4069
rect 28169 4060 28181 4063
rect 27764 4032 28181 4060
rect 27764 4020 27770 4032
rect 28169 4029 28181 4032
rect 28215 4029 28227 4063
rect 28828 4060 28856 4100
rect 28905 4097 28917 4131
rect 28951 4128 28963 4131
rect 29178 4128 29184 4140
rect 28951 4100 29184 4128
rect 28951 4097 28963 4100
rect 28905 4091 28963 4097
rect 29178 4088 29184 4100
rect 29236 4088 29242 4140
rect 29270 4088 29276 4140
rect 29328 4128 29334 4140
rect 29457 4131 29515 4137
rect 29457 4128 29469 4131
rect 29328 4100 29469 4128
rect 29328 4088 29334 4100
rect 29457 4097 29469 4100
rect 29503 4097 29515 4131
rect 29457 4091 29515 4097
rect 29638 4088 29644 4140
rect 29696 4088 29702 4140
rect 30285 4131 30343 4137
rect 30285 4097 30297 4131
rect 30331 4128 30343 4131
rect 30466 4128 30472 4140
rect 30331 4100 30472 4128
rect 30331 4097 30343 4100
rect 30285 4091 30343 4097
rect 30466 4088 30472 4100
rect 30524 4088 30530 4140
rect 30650 4088 30656 4140
rect 30708 4128 30714 4140
rect 30929 4131 30987 4137
rect 30929 4128 30941 4131
rect 30708 4100 30941 4128
rect 30708 4088 30714 4100
rect 30929 4097 30941 4100
rect 30975 4097 30987 4131
rect 30929 4091 30987 4097
rect 32125 4131 32183 4137
rect 32125 4097 32137 4131
rect 32171 4128 32183 4131
rect 32306 4128 32312 4140
rect 32171 4100 32312 4128
rect 32171 4097 32183 4100
rect 32125 4091 32183 4097
rect 32306 4088 32312 4100
rect 32364 4088 32370 4140
rect 32677 4131 32735 4137
rect 32677 4097 32689 4131
rect 32723 4128 32735 4131
rect 33134 4128 33140 4140
rect 32723 4100 33140 4128
rect 32723 4097 32735 4100
rect 32677 4091 32735 4097
rect 33134 4088 33140 4100
rect 33192 4088 33198 4140
rect 33318 4088 33324 4140
rect 33376 4128 33382 4140
rect 33376 4100 37780 4128
rect 33376 4088 33382 4100
rect 29362 4060 29368 4072
rect 28828 4032 29368 4060
rect 28169 4023 28227 4029
rect 29362 4020 29368 4032
rect 29420 4020 29426 4072
rect 30374 4020 30380 4072
rect 30432 4020 30438 4072
rect 31018 4020 31024 4072
rect 31076 4060 31082 4072
rect 31757 4063 31815 4069
rect 31757 4060 31769 4063
rect 31076 4032 31769 4060
rect 31076 4020 31082 4032
rect 31757 4029 31769 4032
rect 31803 4029 31815 4063
rect 31757 4023 31815 4029
rect 32490 4020 32496 4072
rect 32548 4060 32554 4072
rect 33413 4063 33471 4069
rect 33413 4060 33425 4063
rect 32548 4032 33425 4060
rect 32548 4020 32554 4032
rect 33413 4029 33425 4032
rect 33459 4029 33471 4063
rect 33413 4023 33471 4029
rect 33870 4020 33876 4072
rect 33928 4060 33934 4072
rect 34149 4063 34207 4069
rect 34149 4060 34161 4063
rect 33928 4032 34161 4060
rect 33928 4020 33934 4032
rect 34149 4029 34161 4032
rect 34195 4029 34207 4063
rect 34149 4023 34207 4029
rect 34790 4020 34796 4072
rect 34848 4060 34854 4072
rect 34885 4063 34943 4069
rect 34885 4060 34897 4063
rect 34848 4032 34897 4060
rect 34848 4020 34854 4032
rect 34885 4029 34897 4032
rect 34931 4029 34943 4063
rect 34885 4023 34943 4029
rect 34974 4020 34980 4072
rect 35032 4060 35038 4072
rect 35621 4063 35679 4069
rect 35621 4060 35633 4063
rect 35032 4032 35633 4060
rect 35032 4020 35038 4032
rect 35621 4029 35633 4032
rect 35667 4029 35679 4063
rect 35621 4023 35679 4029
rect 35986 4020 35992 4072
rect 36044 4020 36050 4072
rect 37645 4063 37703 4069
rect 37645 4029 37657 4063
rect 37691 4029 37703 4063
rect 37752 4060 37780 4100
rect 37826 4088 37832 4140
rect 37884 4088 37890 4140
rect 38930 4088 38936 4140
rect 38988 4088 38994 4140
rect 43530 4088 43536 4140
rect 43588 4088 43594 4140
rect 44284 4137 44312 4168
rect 46106 4156 46112 4208
rect 46164 4196 46170 4208
rect 55398 4196 55404 4208
rect 46164 4168 55404 4196
rect 46164 4156 46170 4168
rect 55398 4156 55404 4168
rect 55456 4156 55462 4208
rect 55490 4156 55496 4208
rect 55548 4196 55554 4208
rect 68094 4196 68100 4208
rect 55548 4168 68100 4196
rect 55548 4156 55554 4168
rect 68094 4156 68100 4168
rect 68152 4156 68158 4208
rect 44269 4131 44327 4137
rect 44269 4097 44281 4131
rect 44315 4097 44327 4131
rect 44269 4091 44327 4097
rect 47673 4131 47731 4137
rect 47673 4097 47685 4131
rect 47719 4128 47731 4131
rect 47946 4128 47952 4140
rect 47719 4100 47952 4128
rect 47719 4097 47731 4100
rect 47673 4091 47731 4097
rect 47946 4088 47952 4100
rect 48004 4088 48010 4140
rect 48225 4131 48283 4137
rect 48225 4097 48237 4131
rect 48271 4128 48283 4131
rect 53282 4128 53288 4140
rect 48271 4100 53288 4128
rect 48271 4097 48283 4100
rect 48225 4091 48283 4097
rect 53282 4088 53288 4100
rect 53340 4088 53346 4140
rect 53377 4131 53435 4137
rect 53377 4097 53389 4131
rect 53423 4128 53435 4131
rect 55858 4128 55864 4140
rect 53423 4100 55864 4128
rect 53423 4097 53435 4100
rect 53377 4091 53435 4097
rect 55858 4088 55864 4100
rect 55916 4088 55922 4140
rect 38289 4063 38347 4069
rect 38289 4060 38301 4063
rect 37752 4032 38301 4060
rect 37645 4023 37703 4029
rect 38289 4029 38301 4032
rect 38335 4029 38347 4063
rect 38289 4023 38347 4029
rect 42153 4063 42211 4069
rect 42153 4029 42165 4063
rect 42199 4060 42211 4063
rect 42242 4060 42248 4072
rect 42199 4032 42248 4060
rect 42199 4029 42211 4032
rect 42153 4023 42211 4029
rect 37182 3992 37188 4004
rect 27172 3964 37188 3992
rect 37182 3952 37188 3964
rect 37240 3952 37246 4004
rect 37660 3992 37688 4023
rect 42242 4020 42248 4032
rect 42300 4020 42306 4072
rect 42429 4063 42487 4069
rect 42429 4029 42441 4063
rect 42475 4060 42487 4063
rect 43346 4060 43352 4072
rect 42475 4032 43352 4060
rect 42475 4029 42487 4032
rect 42429 4023 42487 4029
rect 43346 4020 43352 4032
rect 43404 4020 43410 4072
rect 45462 4020 45468 4072
rect 45520 4020 45526 4072
rect 47578 4060 47584 4072
rect 46032 4032 47584 4060
rect 41322 3992 41328 4004
rect 37660 3964 41328 3992
rect 41322 3952 41328 3964
rect 41380 3952 41386 4004
rect 44085 3995 44143 4001
rect 44085 3961 44097 3995
rect 44131 3992 44143 3995
rect 46032 3992 46060 4032
rect 47578 4020 47584 4032
rect 47636 4020 47642 4072
rect 47762 4020 47768 4072
rect 47820 4060 47826 4072
rect 49326 4060 49332 4072
rect 47820 4032 49332 4060
rect 47820 4020 47826 4032
rect 49326 4020 49332 4032
rect 49384 4020 49390 4072
rect 49418 4020 49424 4072
rect 49476 4060 49482 4072
rect 52733 4063 52791 4069
rect 52733 4060 52745 4063
rect 49476 4032 52745 4060
rect 49476 4020 49482 4032
rect 52733 4029 52745 4032
rect 52779 4029 52791 4063
rect 52733 4023 52791 4029
rect 44131 3964 46060 3992
rect 46109 3995 46167 4001
rect 44131 3961 44143 3964
rect 44085 3955 44143 3961
rect 46109 3961 46121 3995
rect 46155 3992 46167 3995
rect 51534 3992 51540 4004
rect 46155 3964 51540 3992
rect 46155 3961 46167 3964
rect 46109 3955 46167 3961
rect 51534 3952 51540 3964
rect 51592 3952 51598 4004
rect 52270 3952 52276 4004
rect 52328 3992 52334 4004
rect 58618 3992 58624 4004
rect 52328 3964 58624 3992
rect 52328 3952 52334 3964
rect 58618 3952 58624 3964
rect 58676 3952 58682 4004
rect 25222 3884 25228 3936
rect 25280 3884 25286 3936
rect 25314 3884 25320 3936
rect 25372 3884 25378 3936
rect 26050 3884 26056 3936
rect 26108 3884 26114 3936
rect 28077 3927 28135 3933
rect 28077 3893 28089 3927
rect 28123 3924 28135 3927
rect 28442 3924 28448 3936
rect 28123 3896 28448 3924
rect 28123 3893 28135 3896
rect 28077 3887 28135 3893
rect 28442 3884 28448 3896
rect 28500 3884 28506 3936
rect 28813 3927 28871 3933
rect 28813 3893 28825 3927
rect 28859 3924 28871 3927
rect 28994 3924 29000 3936
rect 28859 3896 29000 3924
rect 28859 3893 28871 3896
rect 28813 3887 28871 3893
rect 28994 3884 29000 3896
rect 29052 3884 29058 3936
rect 29086 3884 29092 3936
rect 29144 3924 29150 3936
rect 30926 3924 30932 3936
rect 29144 3896 30932 3924
rect 29144 3884 29150 3896
rect 30926 3884 30932 3896
rect 30984 3884 30990 3936
rect 31202 3884 31208 3936
rect 31260 3884 31266 3936
rect 32858 3884 32864 3936
rect 32916 3884 32922 3936
rect 33226 3884 33232 3936
rect 33284 3924 33290 3936
rect 33597 3927 33655 3933
rect 33597 3924 33609 3927
rect 33284 3896 33609 3924
rect 33284 3884 33290 3896
rect 33597 3893 33609 3896
rect 33643 3893 33655 3927
rect 33597 3887 33655 3893
rect 34054 3884 34060 3936
rect 34112 3924 34118 3936
rect 34333 3927 34391 3933
rect 34333 3924 34345 3927
rect 34112 3896 34345 3924
rect 34112 3884 34118 3896
rect 34333 3893 34345 3896
rect 34379 3893 34391 3927
rect 34333 3887 34391 3893
rect 35066 3884 35072 3936
rect 35124 3884 35130 3936
rect 36633 3927 36691 3933
rect 36633 3893 36645 3927
rect 36679 3924 36691 3927
rect 36814 3924 36820 3936
rect 36679 3896 36820 3924
rect 36679 3893 36691 3896
rect 36633 3887 36691 3893
rect 36814 3884 36820 3896
rect 36872 3884 36878 3936
rect 41506 3884 41512 3936
rect 41564 3884 41570 3936
rect 42981 3927 43039 3933
rect 42981 3893 42993 3927
rect 43027 3924 43039 3927
rect 43806 3924 43812 3936
rect 43027 3896 43812 3924
rect 43027 3893 43039 3896
rect 42981 3887 43039 3893
rect 43806 3884 43812 3896
rect 43864 3884 43870 3936
rect 44913 3927 44971 3933
rect 44913 3893 44925 3927
rect 44959 3924 44971 3927
rect 50798 3924 50804 3936
rect 44959 3896 50804 3924
rect 44959 3893 44971 3896
rect 44913 3887 44971 3893
rect 50798 3884 50804 3896
rect 50856 3884 50862 3936
rect 55858 3884 55864 3936
rect 55916 3924 55922 3936
rect 65242 3924 65248 3936
rect 55916 3896 65248 3924
rect 55916 3884 55922 3896
rect 65242 3884 65248 3896
rect 65300 3884 65306 3936
rect 1012 3834 74980 3856
rect 1012 3782 1858 3834
rect 1910 3782 1922 3834
rect 1974 3782 1986 3834
rect 2038 3782 2050 3834
rect 2102 3782 2114 3834
rect 2166 3782 11858 3834
rect 11910 3782 11922 3834
rect 11974 3782 11986 3834
rect 12038 3782 12050 3834
rect 12102 3782 12114 3834
rect 12166 3782 21858 3834
rect 21910 3782 21922 3834
rect 21974 3782 21986 3834
rect 22038 3782 22050 3834
rect 22102 3782 22114 3834
rect 22166 3782 31858 3834
rect 31910 3782 31922 3834
rect 31974 3782 31986 3834
rect 32038 3782 32050 3834
rect 32102 3782 32114 3834
rect 32166 3782 41858 3834
rect 41910 3782 41922 3834
rect 41974 3782 41986 3834
rect 42038 3782 42050 3834
rect 42102 3782 42114 3834
rect 42166 3782 51858 3834
rect 51910 3782 51922 3834
rect 51974 3782 51986 3834
rect 52038 3782 52050 3834
rect 52102 3782 52114 3834
rect 52166 3782 61858 3834
rect 61910 3782 61922 3834
rect 61974 3782 61986 3834
rect 62038 3782 62050 3834
rect 62102 3782 62114 3834
rect 62166 3782 71858 3834
rect 71910 3782 71922 3834
rect 71974 3782 71986 3834
rect 72038 3782 72050 3834
rect 72102 3782 72114 3834
rect 72166 3782 74980 3834
rect 1012 3760 74980 3782
rect 27890 3720 27896 3732
rect 25516 3692 27896 3720
rect 23569 3519 23627 3525
rect 23569 3485 23581 3519
rect 23615 3516 23627 3519
rect 23658 3516 23664 3528
rect 23615 3488 23664 3516
rect 23615 3485 23627 3488
rect 23569 3479 23627 3485
rect 23658 3476 23664 3488
rect 23716 3476 23722 3528
rect 24857 3519 24915 3525
rect 24857 3485 24869 3519
rect 24903 3516 24915 3519
rect 25314 3516 25320 3528
rect 24903 3488 25320 3516
rect 24903 3485 24915 3488
rect 24857 3479 24915 3485
rect 25314 3476 25320 3488
rect 25372 3476 25378 3528
rect 25516 3516 25544 3692
rect 27890 3680 27896 3692
rect 27948 3680 27954 3732
rect 29273 3723 29331 3729
rect 29273 3689 29285 3723
rect 29319 3720 29331 3723
rect 29822 3720 29828 3732
rect 29319 3692 29828 3720
rect 29319 3689 29331 3692
rect 29273 3683 29331 3689
rect 29822 3680 29828 3692
rect 29880 3680 29886 3732
rect 29914 3680 29920 3732
rect 29972 3720 29978 3732
rect 30742 3720 30748 3732
rect 29972 3692 30748 3720
rect 29972 3680 29978 3692
rect 30742 3680 30748 3692
rect 30800 3680 30806 3732
rect 31481 3723 31539 3729
rect 31481 3689 31493 3723
rect 31527 3720 31539 3723
rect 33410 3720 33416 3732
rect 31527 3692 33416 3720
rect 31527 3689 31539 3692
rect 31481 3683 31539 3689
rect 33410 3680 33416 3692
rect 33468 3680 33474 3732
rect 35250 3680 35256 3732
rect 35308 3720 35314 3732
rect 35345 3723 35403 3729
rect 35345 3720 35357 3723
rect 35308 3692 35357 3720
rect 35308 3680 35314 3692
rect 35345 3689 35357 3692
rect 35391 3689 35403 3723
rect 40126 3720 40132 3732
rect 35345 3683 35403 3689
rect 35866 3692 40132 3720
rect 29730 3652 29736 3664
rect 27448 3624 29736 3652
rect 25593 3587 25651 3593
rect 25593 3553 25605 3587
rect 25639 3584 25651 3587
rect 27338 3584 27344 3596
rect 25639 3556 27344 3584
rect 25639 3553 25651 3556
rect 25593 3547 25651 3553
rect 27338 3544 27344 3556
rect 27396 3544 27402 3596
rect 25685 3519 25743 3525
rect 25685 3516 25697 3519
rect 25516 3488 25697 3516
rect 25685 3485 25697 3488
rect 25731 3485 25743 3519
rect 25685 3479 25743 3485
rect 26418 3476 26424 3528
rect 26476 3476 26482 3528
rect 27448 3516 27476 3624
rect 29730 3612 29736 3624
rect 29788 3612 29794 3664
rect 35866 3652 35894 3692
rect 40126 3680 40132 3692
rect 40184 3680 40190 3732
rect 40788 3692 42196 3720
rect 29840 3624 35894 3652
rect 27890 3544 27896 3596
rect 27948 3584 27954 3596
rect 29086 3584 29092 3596
rect 27948 3556 29092 3584
rect 27948 3544 27954 3556
rect 29086 3544 29092 3556
rect 29144 3544 29150 3596
rect 29840 3593 29868 3624
rect 29825 3587 29883 3593
rect 29825 3553 29837 3587
rect 29871 3553 29883 3587
rect 32858 3584 32864 3596
rect 29825 3547 29883 3553
rect 30024 3556 32864 3584
rect 26528 3488 27476 3516
rect 24581 3451 24639 3457
rect 24581 3417 24593 3451
rect 24627 3448 24639 3451
rect 26528 3448 26556 3488
rect 27798 3476 27804 3528
rect 27856 3476 27862 3528
rect 27982 3476 27988 3528
rect 28040 3476 28046 3528
rect 30024 3525 30052 3556
rect 32858 3544 32864 3556
rect 32916 3544 32922 3596
rect 34054 3544 34060 3596
rect 34112 3584 34118 3596
rect 34333 3587 34391 3593
rect 34333 3584 34345 3587
rect 34112 3556 34345 3584
rect 34112 3544 34118 3556
rect 34333 3553 34345 3556
rect 34379 3553 34391 3587
rect 34333 3547 34391 3553
rect 38933 3587 38991 3593
rect 38933 3553 38945 3587
rect 38979 3584 38991 3587
rect 40788 3584 40816 3692
rect 40862 3612 40868 3664
rect 40920 3612 40926 3664
rect 42168 3652 42196 3692
rect 42242 3680 42248 3732
rect 42300 3720 42306 3732
rect 42705 3723 42763 3729
rect 42705 3720 42717 3723
rect 42300 3692 42717 3720
rect 42300 3680 42306 3692
rect 42705 3689 42717 3692
rect 42751 3689 42763 3723
rect 42705 3683 42763 3689
rect 43346 3680 43352 3732
rect 43404 3720 43410 3732
rect 43441 3723 43499 3729
rect 43441 3720 43453 3723
rect 43404 3692 43453 3720
rect 43404 3680 43410 3692
rect 43441 3689 43453 3692
rect 43487 3689 43499 3723
rect 48406 3720 48412 3732
rect 43441 3683 43499 3689
rect 46308 3692 48412 3720
rect 45002 3652 45008 3664
rect 42168 3624 45008 3652
rect 45002 3612 45008 3624
rect 45060 3612 45066 3664
rect 38979 3556 40816 3584
rect 38979 3553 38991 3556
rect 38933 3547 38991 3553
rect 41506 3544 41512 3596
rect 41564 3584 41570 3596
rect 41969 3587 42027 3593
rect 41969 3584 41981 3587
rect 41564 3556 41981 3584
rect 41564 3544 41570 3556
rect 41969 3553 41981 3556
rect 42015 3553 42027 3587
rect 41969 3547 42027 3553
rect 42242 3544 42248 3596
rect 42300 3584 42306 3596
rect 43993 3587 44051 3593
rect 43993 3584 44005 3587
rect 42300 3556 44005 3584
rect 42300 3544 42306 3556
rect 43993 3553 44005 3556
rect 44039 3553 44051 3587
rect 43993 3547 44051 3553
rect 44726 3544 44732 3596
rect 44784 3584 44790 3596
rect 45649 3587 45707 3593
rect 45649 3584 45661 3587
rect 44784 3556 45661 3584
rect 44784 3544 44790 3556
rect 45649 3553 45661 3556
rect 45695 3553 45707 3587
rect 45649 3547 45707 3553
rect 28721 3519 28779 3525
rect 28721 3485 28733 3519
rect 28767 3485 28779 3519
rect 28721 3479 28779 3485
rect 30009 3519 30067 3525
rect 30009 3485 30021 3519
rect 30055 3485 30067 3519
rect 30009 3479 30067 3485
rect 30653 3519 30711 3525
rect 30653 3485 30665 3519
rect 30699 3485 30711 3519
rect 30653 3479 30711 3485
rect 30929 3519 30987 3525
rect 30929 3485 30941 3519
rect 30975 3516 30987 3519
rect 32217 3519 32275 3525
rect 30975 3488 32168 3516
rect 30975 3485 30987 3488
rect 30929 3479 30987 3485
rect 24627 3420 26556 3448
rect 24627 3417 24639 3420
rect 24581 3411 24639 3417
rect 26602 3408 26608 3460
rect 26660 3448 26666 3460
rect 27157 3451 27215 3457
rect 27157 3448 27169 3451
rect 26660 3420 27169 3448
rect 26660 3408 26666 3420
rect 27157 3417 27169 3420
rect 27203 3417 27215 3451
rect 28736 3448 28764 3479
rect 30558 3448 30564 3460
rect 28736 3420 30564 3448
rect 27157 3411 27215 3417
rect 30558 3408 30564 3420
rect 30616 3408 30622 3460
rect 24026 3340 24032 3392
rect 24084 3380 24090 3392
rect 24121 3383 24179 3389
rect 24121 3380 24133 3383
rect 24084 3352 24133 3380
rect 24084 3340 24090 3352
rect 24121 3349 24133 3352
rect 24167 3349 24179 3383
rect 24121 3343 24179 3349
rect 24946 3340 24952 3392
rect 25004 3340 25010 3392
rect 26329 3383 26387 3389
rect 26329 3349 26341 3383
rect 26375 3380 26387 3383
rect 26970 3380 26976 3392
rect 26375 3352 26976 3380
rect 26375 3349 26387 3352
rect 26329 3343 26387 3349
rect 26970 3340 26976 3352
rect 27028 3340 27034 3392
rect 27062 3340 27068 3392
rect 27120 3340 27126 3392
rect 28537 3383 28595 3389
rect 28537 3349 28549 3383
rect 28583 3380 28595 3383
rect 29178 3380 29184 3392
rect 28583 3352 29184 3380
rect 28583 3349 28595 3352
rect 28537 3343 28595 3349
rect 29178 3340 29184 3352
rect 29236 3340 29242 3392
rect 30098 3340 30104 3392
rect 30156 3340 30162 3392
rect 30668 3380 30696 3479
rect 30742 3408 30748 3460
rect 30800 3448 30806 3460
rect 31573 3451 31631 3457
rect 31573 3448 31585 3451
rect 30800 3420 31585 3448
rect 30800 3408 30806 3420
rect 31573 3417 31585 3420
rect 31619 3417 31631 3451
rect 31573 3411 31631 3417
rect 31662 3380 31668 3392
rect 30668 3352 31668 3380
rect 31662 3340 31668 3352
rect 31720 3340 31726 3392
rect 32140 3380 32168 3488
rect 32217 3485 32229 3519
rect 32263 3485 32275 3519
rect 32217 3479 32275 3485
rect 32232 3448 32260 3479
rect 32306 3476 32312 3528
rect 32364 3476 32370 3528
rect 32582 3476 32588 3528
rect 32640 3516 32646 3528
rect 33045 3519 33103 3525
rect 33045 3516 33057 3519
rect 32640 3488 33057 3516
rect 32640 3476 32646 3488
rect 33045 3485 33057 3488
rect 33091 3485 33103 3519
rect 33045 3479 33103 3485
rect 34698 3476 34704 3528
rect 34756 3476 34762 3528
rect 35894 3476 35900 3528
rect 35952 3516 35958 3528
rect 35989 3519 36047 3525
rect 35989 3516 36001 3519
rect 35952 3488 36001 3516
rect 35952 3476 35958 3488
rect 35989 3485 36001 3488
rect 36035 3485 36047 3519
rect 35989 3479 36047 3485
rect 36078 3476 36084 3528
rect 36136 3516 36142 3528
rect 36173 3519 36231 3525
rect 36173 3516 36185 3519
rect 36136 3488 36185 3516
rect 36136 3476 36142 3488
rect 36173 3485 36185 3488
rect 36219 3485 36231 3519
rect 36173 3479 36231 3485
rect 36817 3519 36875 3525
rect 36817 3485 36829 3519
rect 36863 3516 36875 3519
rect 37461 3519 37519 3525
rect 37461 3516 37473 3519
rect 36863 3488 37473 3516
rect 36863 3485 36875 3488
rect 36817 3479 36875 3485
rect 37461 3485 37473 3488
rect 37507 3485 37519 3519
rect 37461 3479 37519 3485
rect 38378 3476 38384 3528
rect 38436 3476 38442 3528
rect 39114 3476 39120 3528
rect 39172 3476 39178 3528
rect 40310 3476 40316 3528
rect 40368 3476 40374 3528
rect 40586 3476 40592 3528
rect 40644 3476 40650 3528
rect 41322 3476 41328 3528
rect 41380 3476 41386 3528
rect 41598 3476 41604 3528
rect 41656 3516 41662 3528
rect 43257 3519 43315 3525
rect 43257 3516 43269 3519
rect 41656 3488 43269 3516
rect 41656 3476 41662 3488
rect 43257 3485 43269 3488
rect 43303 3485 43315 3519
rect 43257 3479 43315 3485
rect 44634 3476 44640 3528
rect 44692 3476 44698 3528
rect 45005 3519 45063 3525
rect 45005 3485 45017 3519
rect 45051 3516 45063 3519
rect 45554 3516 45560 3528
rect 45051 3488 45560 3516
rect 45051 3485 45063 3488
rect 45005 3479 45063 3485
rect 45554 3476 45560 3488
rect 45612 3476 45618 3528
rect 46308 3516 46336 3692
rect 48406 3680 48412 3692
rect 48464 3680 48470 3732
rect 49418 3680 49424 3732
rect 49476 3680 49482 3732
rect 49602 3680 49608 3732
rect 49660 3720 49666 3732
rect 55858 3720 55864 3732
rect 49660 3692 55864 3720
rect 49660 3680 49666 3692
rect 55858 3680 55864 3692
rect 55916 3680 55922 3732
rect 65518 3720 65524 3732
rect 55968 3692 65524 3720
rect 48314 3652 48320 3664
rect 46492 3624 48320 3652
rect 46492 3593 46520 3624
rect 48314 3612 48320 3624
rect 48372 3612 48378 3664
rect 54662 3612 54668 3664
rect 54720 3652 54726 3664
rect 55968 3652 55996 3692
rect 65518 3680 65524 3692
rect 65576 3680 65582 3732
rect 54720 3624 55996 3652
rect 54720 3612 54726 3624
rect 59078 3612 59084 3664
rect 59136 3652 59142 3664
rect 63586 3652 63592 3664
rect 59136 3624 63592 3652
rect 59136 3612 59142 3624
rect 63586 3612 63592 3624
rect 63644 3612 63650 3664
rect 64690 3652 64696 3664
rect 64340 3624 64696 3652
rect 46477 3587 46535 3593
rect 46477 3553 46489 3587
rect 46523 3553 46535 3587
rect 46477 3547 46535 3553
rect 47765 3587 47823 3593
rect 47765 3553 47777 3587
rect 47811 3584 47823 3587
rect 49878 3584 49884 3596
rect 47811 3556 49884 3584
rect 47811 3553 47823 3556
rect 47765 3547 47823 3553
rect 49878 3544 49884 3556
rect 49936 3544 49942 3596
rect 50893 3587 50951 3593
rect 50893 3553 50905 3587
rect 50939 3584 50951 3587
rect 53926 3584 53932 3596
rect 50939 3556 53932 3584
rect 50939 3553 50951 3556
rect 50893 3547 50951 3553
rect 53926 3544 53932 3556
rect 53984 3544 53990 3596
rect 64340 3593 64368 3624
rect 64690 3612 64696 3624
rect 64748 3612 64754 3664
rect 64325 3587 64383 3593
rect 64325 3553 64337 3587
rect 64371 3553 64383 3587
rect 64325 3547 64383 3553
rect 46216 3488 46336 3516
rect 47213 3519 47271 3525
rect 33134 3448 33140 3460
rect 32232 3420 33140 3448
rect 33134 3408 33140 3420
rect 33192 3408 33198 3460
rect 35158 3448 35164 3460
rect 33244 3420 35164 3448
rect 32766 3380 32772 3392
rect 32140 3352 32772 3380
rect 32766 3340 32772 3352
rect 32824 3340 32830 3392
rect 32950 3340 32956 3392
rect 33008 3340 33014 3392
rect 33042 3340 33048 3392
rect 33100 3380 33106 3392
rect 33244 3380 33272 3420
rect 35158 3408 35164 3420
rect 35216 3408 35222 3460
rect 35618 3408 35624 3460
rect 35676 3448 35682 3460
rect 36909 3451 36967 3457
rect 36909 3448 36921 3451
rect 35676 3420 36921 3448
rect 35676 3408 35682 3420
rect 36909 3417 36921 3420
rect 36955 3417 36967 3451
rect 36909 3411 36967 3417
rect 41049 3451 41107 3457
rect 41049 3417 41061 3451
rect 41095 3448 41107 3451
rect 42334 3448 42340 3460
rect 41095 3420 42340 3448
rect 41095 3417 41107 3420
rect 41049 3411 41107 3417
rect 42334 3408 42340 3420
rect 42392 3408 42398 3460
rect 44361 3451 44419 3457
rect 44361 3417 44373 3451
rect 44407 3448 44419 3451
rect 46216 3448 46244 3488
rect 47213 3485 47225 3519
rect 47259 3516 47271 3519
rect 47486 3516 47492 3528
rect 47259 3488 47492 3516
rect 47259 3485 47271 3488
rect 47213 3479 47271 3485
rect 47486 3476 47492 3488
rect 47544 3476 47550 3528
rect 47949 3519 48007 3525
rect 47949 3485 47961 3519
rect 47995 3516 48007 3519
rect 48593 3519 48651 3525
rect 48593 3516 48605 3519
rect 47995 3488 48605 3516
rect 47995 3485 48007 3488
rect 47949 3479 48007 3485
rect 48593 3485 48605 3488
rect 48639 3485 48651 3519
rect 48593 3479 48651 3485
rect 48958 3476 48964 3528
rect 49016 3516 49022 3528
rect 49145 3519 49203 3525
rect 49145 3516 49157 3519
rect 49016 3488 49157 3516
rect 49016 3476 49022 3488
rect 49145 3485 49157 3488
rect 49191 3485 49203 3519
rect 49145 3479 49203 3485
rect 49605 3519 49663 3525
rect 49605 3485 49617 3519
rect 49651 3485 49663 3519
rect 49605 3479 49663 3485
rect 44407 3420 46244 3448
rect 46293 3451 46351 3457
rect 44407 3417 44419 3420
rect 44361 3411 44419 3417
rect 46293 3417 46305 3451
rect 46339 3448 46351 3451
rect 47118 3448 47124 3460
rect 46339 3420 47124 3448
rect 46339 3417 46351 3420
rect 46293 3411 46351 3417
rect 47118 3408 47124 3420
rect 47176 3408 47182 3460
rect 49620 3448 49648 3479
rect 50706 3476 50712 3528
rect 50764 3476 50770 3528
rect 51721 3519 51779 3525
rect 51721 3485 51733 3519
rect 51767 3516 51779 3519
rect 52638 3516 52644 3528
rect 51767 3488 52644 3516
rect 51767 3485 51779 3488
rect 51721 3479 51779 3485
rect 52638 3476 52644 3488
rect 52696 3476 52702 3528
rect 53006 3476 53012 3528
rect 53064 3476 53070 3528
rect 55861 3519 55919 3525
rect 55861 3485 55873 3519
rect 55907 3516 55919 3519
rect 55950 3516 55956 3528
rect 55907 3488 55956 3516
rect 55907 3485 55919 3488
rect 55861 3479 55919 3485
rect 55950 3476 55956 3488
rect 56008 3476 56014 3528
rect 57609 3519 57667 3525
rect 57609 3485 57621 3519
rect 57655 3516 57667 3519
rect 60366 3516 60372 3528
rect 57655 3488 60372 3516
rect 57655 3485 57667 3488
rect 57609 3479 57667 3485
rect 60366 3476 60372 3488
rect 60424 3476 60430 3528
rect 60461 3519 60519 3525
rect 60461 3485 60473 3519
rect 60507 3516 60519 3519
rect 64509 3519 64567 3525
rect 60507 3488 64460 3516
rect 60507 3485 60519 3488
rect 60461 3479 60519 3485
rect 51534 3448 51540 3460
rect 49620 3420 51540 3448
rect 51534 3408 51540 3420
rect 51592 3408 51598 3460
rect 52273 3451 52331 3457
rect 52273 3417 52285 3451
rect 52319 3448 52331 3451
rect 54018 3448 54024 3460
rect 52319 3420 54024 3448
rect 52319 3417 52331 3420
rect 52273 3411 52331 3417
rect 54018 3408 54024 3420
rect 54076 3408 54082 3460
rect 58621 3451 58679 3457
rect 58621 3417 58633 3451
rect 58667 3448 58679 3451
rect 59170 3448 59176 3460
rect 58667 3420 59176 3448
rect 58667 3417 58679 3420
rect 58621 3411 58679 3417
rect 59170 3408 59176 3420
rect 59228 3408 59234 3460
rect 60476 3420 60688 3448
rect 33100 3352 33272 3380
rect 33100 3340 33106 3352
rect 33686 3340 33692 3392
rect 33744 3340 33750 3392
rect 33778 3340 33784 3392
rect 33836 3340 33842 3392
rect 34882 3340 34888 3392
rect 34940 3380 34946 3392
rect 35437 3383 35495 3389
rect 35437 3380 35449 3383
rect 34940 3352 35449 3380
rect 34940 3340 34946 3352
rect 35437 3349 35449 3352
rect 35483 3349 35495 3383
rect 35437 3343 35495 3349
rect 37458 3340 37464 3392
rect 37516 3380 37522 3392
rect 37829 3383 37887 3389
rect 37829 3380 37841 3383
rect 37516 3352 37841 3380
rect 37516 3340 37522 3352
rect 37829 3349 37841 3352
rect 37875 3349 37887 3383
rect 37829 3343 37887 3349
rect 41877 3383 41935 3389
rect 41877 3349 41889 3383
rect 41923 3380 41935 3383
rect 42518 3380 42524 3392
rect 41923 3352 42524 3380
rect 41923 3349 41935 3352
rect 41877 3343 41935 3349
rect 42518 3340 42524 3352
rect 42576 3340 42582 3392
rect 42613 3383 42671 3389
rect 42613 3349 42625 3383
rect 42659 3380 42671 3383
rect 43438 3380 43444 3392
rect 42659 3352 43444 3380
rect 42659 3349 42671 3352
rect 42613 3343 42671 3349
rect 43438 3340 43444 3352
rect 43496 3340 43502 3392
rect 43530 3340 43536 3392
rect 43588 3380 43594 3392
rect 45462 3380 45468 3392
rect 43588 3352 45468 3380
rect 43588 3340 43594 3352
rect 45462 3340 45468 3352
rect 45520 3340 45526 3392
rect 45557 3383 45615 3389
rect 45557 3349 45569 3383
rect 45603 3380 45615 3383
rect 46934 3380 46940 3392
rect 45603 3352 46940 3380
rect 45603 3349 45615 3352
rect 45557 3343 45615 3349
rect 46934 3340 46940 3352
rect 46992 3340 46998 3392
rect 47026 3340 47032 3392
rect 47084 3340 47090 3392
rect 48501 3383 48559 3389
rect 48501 3349 48513 3383
rect 48547 3380 48559 3383
rect 49970 3380 49976 3392
rect 48547 3352 49976 3380
rect 48547 3349 48559 3352
rect 48501 3343 48559 3349
rect 49970 3340 49976 3352
rect 50028 3340 50034 3392
rect 50065 3383 50123 3389
rect 50065 3349 50077 3383
rect 50111 3380 50123 3383
rect 50430 3380 50436 3392
rect 50111 3352 50436 3380
rect 50111 3349 50123 3352
rect 50065 3343 50123 3349
rect 50430 3340 50436 3352
rect 50488 3340 50494 3392
rect 51442 3340 51448 3392
rect 51500 3340 51506 3392
rect 52362 3340 52368 3392
rect 52420 3340 52426 3392
rect 55217 3383 55275 3389
rect 55217 3349 55229 3383
rect 55263 3380 55275 3383
rect 55582 3380 55588 3392
rect 55263 3352 55588 3380
rect 55263 3349 55275 3352
rect 55217 3343 55275 3349
rect 55582 3340 55588 3352
rect 55640 3340 55646 3392
rect 58158 3340 58164 3392
rect 58216 3340 58222 3392
rect 58529 3383 58587 3389
rect 58529 3349 58541 3383
rect 58575 3380 58587 3383
rect 60476 3380 60504 3420
rect 58575 3352 60504 3380
rect 60660 3380 60688 3420
rect 60734 3408 60740 3460
rect 60792 3448 60798 3460
rect 60829 3451 60887 3457
rect 60829 3448 60841 3451
rect 60792 3420 60841 3448
rect 60792 3408 60798 3420
rect 60829 3417 60841 3420
rect 60875 3417 60887 3451
rect 64432 3448 64460 3488
rect 64509 3485 64521 3519
rect 64555 3516 64567 3519
rect 64690 3516 64696 3528
rect 64555 3488 64696 3516
rect 64555 3485 64567 3488
rect 64509 3479 64567 3485
rect 64690 3476 64696 3488
rect 64748 3476 64754 3528
rect 64966 3476 64972 3528
rect 65024 3516 65030 3528
rect 72418 3516 72424 3528
rect 65024 3488 72424 3516
rect 65024 3476 65030 3488
rect 72418 3476 72424 3488
rect 72476 3476 72482 3528
rect 70578 3448 70584 3460
rect 64432 3420 70584 3448
rect 60829 3411 60887 3417
rect 70578 3408 70584 3420
rect 70636 3408 70642 3460
rect 72510 3380 72516 3392
rect 60660 3352 72516 3380
rect 58575 3349 58587 3352
rect 58529 3343 58587 3349
rect 72510 3340 72516 3352
rect 72568 3340 72574 3392
rect 1012 3290 74980 3312
rect 1012 3238 4210 3290
rect 4262 3238 4274 3290
rect 4326 3238 4338 3290
rect 4390 3238 4402 3290
rect 4454 3238 4466 3290
rect 4518 3238 14210 3290
rect 14262 3238 14274 3290
rect 14326 3238 14338 3290
rect 14390 3238 14402 3290
rect 14454 3238 14466 3290
rect 14518 3238 24210 3290
rect 24262 3238 24274 3290
rect 24326 3238 24338 3290
rect 24390 3238 24402 3290
rect 24454 3238 24466 3290
rect 24518 3238 34210 3290
rect 34262 3238 34274 3290
rect 34326 3238 34338 3290
rect 34390 3238 34402 3290
rect 34454 3238 34466 3290
rect 34518 3238 44210 3290
rect 44262 3238 44274 3290
rect 44326 3238 44338 3290
rect 44390 3238 44402 3290
rect 44454 3238 44466 3290
rect 44518 3238 54210 3290
rect 54262 3238 54274 3290
rect 54326 3238 54338 3290
rect 54390 3238 54402 3290
rect 54454 3238 54466 3290
rect 54518 3238 64210 3290
rect 64262 3238 64274 3290
rect 64326 3238 64338 3290
rect 64390 3238 64402 3290
rect 64454 3238 64466 3290
rect 64518 3238 74210 3290
rect 74262 3238 74274 3290
rect 74326 3238 74338 3290
rect 74390 3238 74402 3290
rect 74454 3238 74466 3290
rect 74518 3238 74980 3290
rect 1012 3216 74980 3238
rect 23017 3179 23075 3185
rect 23017 3145 23029 3179
rect 23063 3176 23075 3179
rect 24578 3176 24584 3188
rect 23063 3148 24584 3176
rect 23063 3145 23075 3148
rect 23017 3139 23075 3145
rect 24578 3136 24584 3148
rect 24636 3136 24642 3188
rect 27062 3136 27068 3188
rect 27120 3176 27126 3188
rect 31849 3179 31907 3185
rect 27120 3148 29776 3176
rect 27120 3136 27126 3148
rect 24489 3111 24547 3117
rect 24489 3077 24501 3111
rect 24535 3108 24547 3111
rect 25958 3108 25964 3120
rect 24535 3080 25964 3108
rect 24535 3077 24547 3080
rect 24489 3071 24547 3077
rect 25958 3068 25964 3080
rect 26016 3068 26022 3120
rect 27614 3068 27620 3120
rect 27672 3108 27678 3120
rect 27672 3080 28106 3108
rect 27672 3068 27678 3080
rect 29178 3068 29184 3120
rect 29236 3108 29242 3120
rect 29273 3111 29331 3117
rect 29273 3108 29285 3111
rect 29236 3080 29285 3108
rect 29236 3068 29242 3080
rect 29273 3077 29285 3080
rect 29319 3077 29331 3111
rect 29273 3071 29331 3077
rect 23753 3043 23811 3049
rect 23753 3009 23765 3043
rect 23799 3040 23811 3043
rect 25038 3040 25044 3052
rect 23799 3012 25044 3040
rect 23799 3009 23811 3012
rect 23753 3003 23811 3009
rect 25038 3000 25044 3012
rect 25096 3000 25102 3052
rect 29748 3049 29776 3148
rect 31849 3145 31861 3179
rect 31895 3176 31907 3179
rect 32214 3176 32220 3188
rect 31895 3148 32220 3176
rect 31895 3145 31907 3148
rect 31849 3139 31907 3145
rect 32214 3136 32220 3148
rect 32272 3136 32278 3188
rect 32490 3176 32496 3188
rect 32324 3148 32496 3176
rect 31113 3111 31171 3117
rect 31113 3077 31125 3111
rect 31159 3108 31171 3111
rect 32324 3108 32352 3148
rect 32490 3136 32496 3148
rect 32548 3136 32554 3188
rect 32582 3136 32588 3188
rect 32640 3136 32646 3188
rect 34701 3179 34759 3185
rect 34701 3145 34713 3179
rect 34747 3176 34759 3179
rect 34974 3176 34980 3188
rect 34747 3148 34980 3176
rect 34747 3145 34759 3148
rect 34701 3139 34759 3145
rect 34974 3136 34980 3148
rect 35032 3136 35038 3188
rect 35437 3179 35495 3185
rect 35437 3145 35449 3179
rect 35483 3176 35495 3179
rect 35986 3176 35992 3188
rect 35483 3148 35992 3176
rect 35483 3145 35495 3148
rect 35437 3139 35495 3145
rect 35986 3136 35992 3148
rect 36044 3136 36050 3188
rect 36265 3179 36323 3185
rect 36265 3145 36277 3179
rect 36311 3176 36323 3179
rect 36354 3176 36360 3188
rect 36311 3148 36360 3176
rect 36311 3145 36323 3148
rect 36265 3139 36323 3145
rect 36354 3136 36360 3148
rect 36412 3136 36418 3188
rect 38010 3136 38016 3188
rect 38068 3136 38074 3188
rect 39761 3179 39819 3185
rect 39761 3145 39773 3179
rect 39807 3176 39819 3179
rect 39807 3148 42288 3176
rect 39807 3145 39819 3148
rect 39761 3139 39819 3145
rect 31159 3080 32352 3108
rect 32401 3111 32459 3117
rect 31159 3077 31171 3080
rect 31113 3071 31171 3077
rect 32401 3077 32413 3111
rect 32447 3108 32459 3111
rect 33321 3111 33379 3117
rect 33321 3108 33333 3111
rect 32447 3080 33333 3108
rect 32447 3077 32459 3080
rect 32401 3071 32459 3077
rect 33321 3077 33333 3080
rect 33367 3077 33379 3111
rect 40218 3108 40224 3120
rect 33321 3071 33379 3077
rect 33980 3080 40224 3108
rect 25225 3043 25283 3049
rect 25225 3009 25237 3043
rect 25271 3040 25283 3043
rect 26697 3043 26755 3049
rect 25271 3012 26234 3040
rect 25271 3009 25283 3012
rect 25225 3003 25283 3009
rect 22370 2932 22376 2984
rect 22428 2932 22434 2984
rect 23106 2932 23112 2984
rect 23164 2932 23170 2984
rect 23842 2932 23848 2984
rect 23900 2932 23906 2984
rect 25314 2932 25320 2984
rect 25372 2932 25378 2984
rect 26206 2972 26234 3012
rect 26697 3009 26709 3043
rect 26743 3040 26755 3043
rect 29733 3043 29791 3049
rect 26743 3012 28120 3040
rect 26743 3009 26755 3012
rect 26697 3003 26755 3009
rect 26206 2944 27108 2972
rect 20990 2864 20996 2916
rect 21048 2904 21054 2916
rect 23566 2904 23572 2916
rect 21048 2876 23572 2904
rect 21048 2864 21054 2876
rect 23566 2864 23572 2876
rect 23624 2864 23630 2916
rect 25961 2907 26019 2913
rect 25961 2873 25973 2907
rect 26007 2904 26019 2907
rect 27080 2904 27108 2944
rect 27154 2932 27160 2984
rect 27212 2932 27218 2984
rect 27709 2975 27767 2981
rect 27709 2941 27721 2975
rect 27755 2972 27767 2975
rect 27890 2972 27896 2984
rect 27755 2944 27896 2972
rect 27755 2941 27767 2944
rect 27709 2935 27767 2941
rect 27890 2932 27896 2944
rect 27948 2932 27954 2984
rect 28092 2972 28120 3012
rect 29733 3009 29745 3043
rect 29779 3009 29791 3043
rect 29733 3003 29791 3009
rect 29822 3000 29828 3052
rect 29880 3040 29886 3052
rect 29880 3012 30604 3040
rect 29880 3000 29886 3012
rect 29270 2972 29276 2984
rect 28092 2944 29276 2972
rect 29270 2932 29276 2944
rect 29328 2932 29334 2984
rect 29549 2975 29607 2981
rect 29549 2941 29561 2975
rect 29595 2941 29607 2975
rect 29549 2935 29607 2941
rect 28166 2904 28172 2916
rect 26007 2876 26234 2904
rect 27080 2876 28172 2904
rect 26007 2873 26019 2876
rect 25961 2867 26019 2873
rect 22278 2796 22284 2848
rect 22336 2836 22342 2848
rect 23474 2836 23480 2848
rect 22336 2808 23480 2836
rect 22336 2796 22342 2808
rect 23474 2796 23480 2808
rect 23532 2796 23538 2848
rect 24578 2796 24584 2848
rect 24636 2796 24642 2848
rect 25406 2796 25412 2848
rect 25464 2836 25470 2848
rect 26053 2839 26111 2845
rect 26053 2836 26065 2839
rect 25464 2808 26065 2836
rect 25464 2796 25470 2808
rect 26053 2805 26065 2808
rect 26099 2805 26111 2839
rect 26206 2836 26234 2876
rect 28166 2864 28172 2876
rect 28224 2864 28230 2916
rect 29564 2904 29592 2935
rect 30466 2932 30472 2984
rect 30524 2932 30530 2984
rect 30576 2972 30604 3012
rect 31202 3000 31208 3052
rect 31260 3000 31266 3052
rect 33042 3040 33048 3052
rect 31312 3012 33048 3040
rect 31312 2972 31340 3012
rect 33042 3000 33048 3012
rect 33100 3000 33106 3052
rect 33226 3000 33232 3052
rect 33284 3000 33290 3052
rect 33686 3000 33692 3052
rect 33744 3040 33750 3052
rect 33873 3043 33931 3049
rect 33873 3040 33885 3043
rect 33744 3012 33885 3040
rect 33744 3000 33750 3012
rect 33873 3009 33885 3012
rect 33919 3009 33931 3043
rect 33873 3003 33931 3009
rect 30576 2944 31340 2972
rect 32125 2975 32183 2981
rect 32125 2941 32137 2975
rect 32171 2972 32183 2975
rect 33980 2972 34008 3080
rect 40218 3068 40224 3080
rect 40276 3068 40282 3120
rect 42260 3108 42288 3148
rect 42334 3136 42340 3188
rect 42392 3136 42398 3188
rect 44634 3136 44640 3188
rect 44692 3176 44698 3188
rect 45281 3179 45339 3185
rect 45281 3176 45293 3179
rect 44692 3148 45293 3176
rect 44692 3136 44698 3148
rect 45281 3145 45293 3148
rect 45327 3145 45339 3179
rect 45281 3139 45339 3145
rect 46845 3179 46903 3185
rect 46845 3145 46857 3179
rect 46891 3145 46903 3179
rect 46845 3139 46903 3145
rect 43530 3108 43536 3120
rect 42260 3080 43536 3108
rect 43530 3068 43536 3080
rect 43588 3068 43594 3120
rect 46860 3108 46888 3139
rect 47486 3136 47492 3188
rect 47544 3136 47550 3188
rect 48958 3136 48964 3188
rect 49016 3136 49022 3188
rect 52181 3179 52239 3185
rect 52181 3145 52193 3179
rect 52227 3176 52239 3179
rect 52227 3148 52592 3176
rect 52227 3145 52239 3148
rect 52181 3139 52239 3145
rect 51350 3108 51356 3120
rect 46860 3080 51356 3108
rect 51350 3068 51356 3080
rect 51408 3068 51414 3120
rect 52273 3111 52331 3117
rect 52273 3077 52285 3111
rect 52319 3108 52331 3111
rect 52362 3108 52368 3120
rect 52319 3080 52368 3108
rect 52319 3077 52331 3080
rect 52273 3071 52331 3077
rect 52362 3068 52368 3080
rect 52420 3068 52426 3120
rect 52564 3108 52592 3148
rect 52638 3136 52644 3188
rect 52696 3136 52702 3188
rect 57333 3179 57391 3185
rect 57333 3145 57345 3179
rect 57379 3176 57391 3179
rect 57379 3148 59400 3176
rect 57379 3145 57391 3148
rect 57333 3139 57391 3145
rect 53834 3108 53840 3120
rect 52564 3080 53840 3108
rect 53834 3068 53840 3080
rect 53892 3068 53898 3120
rect 57425 3111 57483 3117
rect 57425 3077 57437 3111
rect 57471 3108 57483 3111
rect 59262 3108 59268 3120
rect 57471 3080 59268 3108
rect 57471 3077 57483 3080
rect 57425 3071 57483 3077
rect 59262 3068 59268 3080
rect 59320 3068 59326 3120
rect 34882 3000 34888 3052
rect 34940 3000 34946 3052
rect 35618 3000 35624 3052
rect 35676 3000 35682 3052
rect 36814 3000 36820 3052
rect 36872 3000 36878 3052
rect 39850 3000 39856 3052
rect 39908 3000 39914 3052
rect 40034 3000 40040 3052
rect 40092 3040 40098 3052
rect 40865 3043 40923 3049
rect 40865 3040 40877 3043
rect 40092 3012 40877 3040
rect 40092 3000 40098 3012
rect 40865 3009 40877 3012
rect 40911 3009 40923 3043
rect 40865 3003 40923 3009
rect 42061 3043 42119 3049
rect 42061 3009 42073 3043
rect 42107 3009 42119 3043
rect 42061 3003 42119 3009
rect 32171 2944 34008 2972
rect 34149 2975 34207 2981
rect 32171 2941 32183 2944
rect 32125 2935 32183 2941
rect 34149 2941 34161 2975
rect 34195 2972 34207 2975
rect 34974 2972 34980 2984
rect 34195 2944 34980 2972
rect 34195 2941 34207 2944
rect 34149 2935 34207 2941
rect 34974 2932 34980 2944
rect 35032 2932 35038 2984
rect 37274 2932 37280 2984
rect 37332 2932 37338 2984
rect 37921 2975 37979 2981
rect 37921 2941 37933 2975
rect 37967 2972 37979 2975
rect 38565 2975 38623 2981
rect 38565 2972 38577 2975
rect 37967 2944 38577 2972
rect 37967 2941 37979 2944
rect 37921 2935 37979 2941
rect 38565 2941 38577 2944
rect 38611 2941 38623 2975
rect 38565 2935 38623 2941
rect 39393 2975 39451 2981
rect 39393 2941 39405 2975
rect 39439 2972 39451 2975
rect 40126 2972 40132 2984
rect 39439 2944 40132 2972
rect 39439 2941 39451 2944
rect 39393 2935 39451 2941
rect 40126 2932 40132 2944
rect 40184 2932 40190 2984
rect 40218 2932 40224 2984
rect 40276 2932 40282 2984
rect 41690 2904 41696 2916
rect 29564 2876 41696 2904
rect 41690 2864 41696 2876
rect 41748 2864 41754 2916
rect 42076 2904 42104 3003
rect 43806 3000 43812 3052
rect 43864 3000 43870 3052
rect 47029 3043 47087 3049
rect 47029 3009 47041 3043
rect 47075 3040 47087 3043
rect 48225 3043 48283 3049
rect 48225 3040 48237 3043
rect 47075 3012 48237 3040
rect 47075 3009 47087 3012
rect 47029 3003 47087 3009
rect 48225 3009 48237 3012
rect 48271 3009 48283 3043
rect 48225 3003 48283 3009
rect 48866 3000 48872 3052
rect 48924 3040 48930 3052
rect 49697 3043 49755 3049
rect 49697 3040 49709 3043
rect 48924 3012 49709 3040
rect 48924 3000 48930 3012
rect 49697 3009 49709 3012
rect 49743 3009 49755 3043
rect 49697 3003 49755 3009
rect 50430 3000 50436 3052
rect 50488 3000 50494 3052
rect 51718 3000 51724 3052
rect 51776 3040 51782 3052
rect 53193 3043 53251 3049
rect 53193 3040 53205 3043
rect 51776 3012 53205 3040
rect 51776 3000 51782 3012
rect 53193 3009 53205 3012
rect 53239 3009 53251 3043
rect 53193 3003 53251 3009
rect 53469 3043 53527 3049
rect 53469 3009 53481 3043
rect 53515 3040 53527 3043
rect 54938 3040 54944 3052
rect 53515 3012 54944 3040
rect 53515 3009 53527 3012
rect 53469 3003 53527 3009
rect 54938 3000 54944 3012
rect 54996 3000 55002 3052
rect 55582 3000 55588 3052
rect 55640 3000 55646 3052
rect 58158 3000 58164 3052
rect 58216 3040 58222 3052
rect 58529 3043 58587 3049
rect 58529 3040 58541 3043
rect 58216 3012 58541 3040
rect 58216 3000 58222 3012
rect 58529 3009 58541 3012
rect 58575 3009 58587 3043
rect 58529 3003 58587 3009
rect 59170 3000 59176 3052
rect 59228 3000 59234 3052
rect 59372 3040 59400 3148
rect 60734 3136 60740 3188
rect 60792 3136 60798 3188
rect 70946 3176 70952 3188
rect 61488 3148 70952 3176
rect 61488 3040 61516 3148
rect 70946 3136 70952 3148
rect 71004 3136 71010 3188
rect 62209 3111 62267 3117
rect 62209 3077 62221 3111
rect 62255 3108 62267 3111
rect 64966 3108 64972 3120
rect 62255 3080 64972 3108
rect 62255 3077 62267 3080
rect 62209 3071 62267 3077
rect 64966 3068 64972 3080
rect 65024 3068 65030 3120
rect 68281 3111 68339 3117
rect 68281 3077 68293 3111
rect 68327 3108 68339 3111
rect 68370 3108 68376 3120
rect 68327 3080 68376 3108
rect 68327 3077 68339 3080
rect 68281 3071 68339 3077
rect 68370 3068 68376 3080
rect 68428 3068 68434 3120
rect 59372 3012 61516 3040
rect 62577 3043 62635 3049
rect 62577 3009 62589 3043
rect 62623 3040 62635 3043
rect 63402 3040 63408 3052
rect 62623 3012 63408 3040
rect 62623 3009 62635 3012
rect 62577 3003 62635 3009
rect 63402 3000 63408 3012
rect 63460 3000 63466 3052
rect 64509 3043 64567 3049
rect 64509 3009 64521 3043
rect 64555 3040 64567 3043
rect 66806 3040 66812 3052
rect 64555 3012 66812 3040
rect 64555 3009 64567 3012
rect 64509 3003 64567 3009
rect 66806 3000 66812 3012
rect 66864 3000 66870 3052
rect 68557 3043 68615 3049
rect 68557 3009 68569 3043
rect 68603 3040 68615 3043
rect 69106 3040 69112 3052
rect 68603 3012 69112 3040
rect 68603 3009 68615 3012
rect 68557 3003 68615 3009
rect 69106 3000 69112 3012
rect 69164 3000 69170 3052
rect 69569 3043 69627 3049
rect 69569 3009 69581 3043
rect 69615 3040 69627 3043
rect 72694 3040 72700 3052
rect 69615 3012 72700 3040
rect 69615 3009 69627 3012
rect 69569 3003 69627 3009
rect 72694 3000 72700 3012
rect 72752 3000 72758 3052
rect 42978 2932 42984 2984
rect 43036 2932 43042 2984
rect 43717 2975 43775 2981
rect 43717 2941 43729 2975
rect 43763 2941 43775 2975
rect 43717 2935 43775 2941
rect 43073 2907 43131 2913
rect 43073 2904 43085 2907
rect 42076 2876 43085 2904
rect 43073 2873 43085 2876
rect 43119 2873 43131 2907
rect 43732 2904 43760 2935
rect 44634 2932 44640 2984
rect 44692 2932 44698 2984
rect 45189 2975 45247 2981
rect 45189 2941 45201 2975
rect 45235 2972 45247 2975
rect 45833 2975 45891 2981
rect 45833 2972 45845 2975
rect 45235 2944 45845 2972
rect 45235 2941 45247 2944
rect 45189 2935 45247 2941
rect 45833 2941 45845 2944
rect 45879 2941 45891 2975
rect 45833 2935 45891 2941
rect 46106 2932 46112 2984
rect 46164 2932 46170 2984
rect 46661 2975 46719 2981
rect 46661 2941 46673 2975
rect 46707 2972 46719 2975
rect 46842 2972 46848 2984
rect 46707 2944 46848 2972
rect 46707 2941 46719 2944
rect 46661 2935 46719 2941
rect 46842 2932 46848 2944
rect 46900 2932 46906 2984
rect 48041 2975 48099 2981
rect 48041 2941 48053 2975
rect 48087 2941 48099 2975
rect 48041 2935 48099 2941
rect 45370 2904 45376 2916
rect 43732 2876 45376 2904
rect 43073 2867 43131 2873
rect 45370 2864 45376 2876
rect 45428 2864 45434 2916
rect 46014 2864 46020 2916
rect 46072 2904 46078 2916
rect 48056 2904 48084 2935
rect 48774 2932 48780 2984
rect 48832 2932 48838 2984
rect 49326 2932 49332 2984
rect 49384 2972 49390 2984
rect 49513 2975 49571 2981
rect 49513 2972 49525 2975
rect 49384 2944 49525 2972
rect 49384 2932 49390 2944
rect 49513 2941 49525 2944
rect 49559 2941 49571 2975
rect 51626 2972 51632 2984
rect 49513 2935 49571 2941
rect 49620 2944 51632 2972
rect 46072 2876 48084 2904
rect 46072 2864 46078 2876
rect 27522 2836 27528 2848
rect 26206 2808 27528 2836
rect 26053 2799 26111 2805
rect 27522 2796 27528 2808
rect 27580 2796 27586 2848
rect 27801 2839 27859 2845
rect 27801 2805 27813 2839
rect 27847 2836 27859 2839
rect 28074 2836 28080 2848
rect 27847 2808 28080 2836
rect 27847 2805 27859 2808
rect 27801 2799 27859 2805
rect 28074 2796 28080 2808
rect 28132 2836 28138 2848
rect 30006 2836 30012 2848
rect 28132 2808 30012 2836
rect 28132 2796 28138 2808
rect 30006 2796 30012 2808
rect 30064 2796 30070 2848
rect 30377 2839 30435 2845
rect 30377 2805 30389 2839
rect 30423 2836 30435 2839
rect 33962 2836 33968 2848
rect 30423 2808 33968 2836
rect 30423 2805 30435 2808
rect 30377 2799 30435 2805
rect 33962 2796 33968 2808
rect 34020 2796 34026 2848
rect 36170 2796 36176 2848
rect 36228 2796 36234 2848
rect 38746 2796 38752 2848
rect 38804 2796 38810 2848
rect 40773 2839 40831 2845
rect 40773 2805 40785 2839
rect 40819 2836 40831 2839
rect 41414 2836 41420 2848
rect 40819 2808 41420 2836
rect 40819 2805 40831 2808
rect 40773 2799 40831 2805
rect 41414 2796 41420 2808
rect 41472 2796 41478 2848
rect 41506 2796 41512 2848
rect 41564 2796 41570 2848
rect 41969 2839 42027 2845
rect 41969 2805 41981 2839
rect 42015 2836 42027 2839
rect 42334 2836 42340 2848
rect 42015 2808 42340 2836
rect 42015 2805 42027 2808
rect 41969 2799 42027 2805
rect 42334 2796 42340 2808
rect 42392 2796 42398 2848
rect 44453 2839 44511 2845
rect 44453 2805 44465 2839
rect 44499 2836 44511 2839
rect 45922 2836 45928 2848
rect 44499 2808 45928 2836
rect 44499 2805 44511 2808
rect 44453 2799 44511 2805
rect 45922 2796 45928 2808
rect 45980 2796 45986 2848
rect 47394 2796 47400 2848
rect 47452 2836 47458 2848
rect 49620 2836 49648 2944
rect 51626 2932 51632 2944
rect 51684 2932 51690 2984
rect 51813 2975 51871 2981
rect 51813 2941 51825 2975
rect 51859 2972 51871 2975
rect 52638 2972 52644 2984
rect 51859 2944 52644 2972
rect 51859 2941 51871 2944
rect 51813 2935 51871 2941
rect 52638 2932 52644 2944
rect 52696 2932 52702 2984
rect 54021 2975 54079 2981
rect 54021 2941 54033 2975
rect 54067 2972 54079 2975
rect 54113 2975 54171 2981
rect 54113 2972 54125 2975
rect 54067 2944 54125 2972
rect 54067 2941 54079 2944
rect 54021 2935 54079 2941
rect 54113 2941 54125 2944
rect 54159 2941 54171 2975
rect 54113 2935 54171 2941
rect 54570 2932 54576 2984
rect 54628 2972 54634 2984
rect 54849 2975 54907 2981
rect 54849 2972 54861 2975
rect 54628 2944 54861 2972
rect 54628 2932 54634 2944
rect 54849 2941 54861 2944
rect 54895 2941 54907 2975
rect 54849 2935 54907 2941
rect 55674 2932 55680 2984
rect 55732 2972 55738 2984
rect 56321 2975 56379 2981
rect 56321 2972 56333 2975
rect 55732 2944 56333 2972
rect 55732 2932 55738 2944
rect 56321 2941 56333 2944
rect 56367 2941 56379 2975
rect 56321 2935 56379 2941
rect 57054 2932 57060 2984
rect 57112 2972 57118 2984
rect 57793 2975 57851 2981
rect 57793 2972 57805 2975
rect 57112 2944 57805 2972
rect 57112 2932 57118 2944
rect 57793 2941 57805 2944
rect 57839 2941 57851 2975
rect 59265 2975 59323 2981
rect 59265 2972 59277 2975
rect 57793 2935 57851 2941
rect 58544 2944 59277 2972
rect 58544 2916 58572 2944
rect 59265 2941 59277 2944
rect 59311 2941 59323 2975
rect 59265 2935 59323 2941
rect 59814 2932 59820 2984
rect 59872 2972 59878 2984
rect 60001 2975 60059 2981
rect 60001 2972 60013 2975
rect 59872 2944 60013 2972
rect 59872 2932 59878 2944
rect 60001 2941 60013 2944
rect 60047 2941 60059 2975
rect 60001 2935 60059 2941
rect 61378 2932 61384 2984
rect 61436 2932 61442 2984
rect 61562 2932 61568 2984
rect 61620 2932 61626 2984
rect 63221 2975 63279 2981
rect 63221 2941 63233 2975
rect 63267 2972 63279 2975
rect 63310 2972 63316 2984
rect 63267 2944 63316 2972
rect 63267 2941 63279 2944
rect 63221 2935 63279 2941
rect 63310 2932 63316 2944
rect 63368 2932 63374 2984
rect 63773 2975 63831 2981
rect 63773 2941 63785 2975
rect 63819 2972 63831 2975
rect 63865 2975 63923 2981
rect 63865 2972 63877 2975
rect 63819 2944 63877 2972
rect 63819 2941 63831 2944
rect 63773 2935 63831 2941
rect 63865 2941 63877 2944
rect 63911 2941 63923 2975
rect 63865 2935 63923 2941
rect 65242 2932 65248 2984
rect 65300 2932 65306 2984
rect 65705 2975 65763 2981
rect 65705 2941 65717 2975
rect 65751 2941 65763 2975
rect 65705 2935 65763 2941
rect 66257 2975 66315 2981
rect 66257 2941 66269 2975
rect 66303 2972 66315 2975
rect 66349 2975 66407 2981
rect 66349 2972 66361 2975
rect 66303 2944 66361 2972
rect 66303 2941 66315 2944
rect 66257 2935 66315 2941
rect 66349 2941 66361 2944
rect 66395 2941 66407 2975
rect 66349 2935 66407 2941
rect 67177 2975 67235 2981
rect 67177 2941 67189 2975
rect 67223 2941 67235 2975
rect 67177 2935 67235 2941
rect 50341 2907 50399 2913
rect 50341 2873 50353 2907
rect 50387 2904 50399 2907
rect 51350 2904 51356 2916
rect 50387 2876 51356 2904
rect 50387 2873 50399 2876
rect 50341 2867 50399 2873
rect 51350 2864 51356 2876
rect 51408 2864 51414 2916
rect 52914 2864 52920 2916
rect 52972 2904 52978 2916
rect 55306 2904 55312 2916
rect 52972 2876 55312 2904
rect 52972 2864 52978 2876
rect 55306 2864 55312 2876
rect 55364 2864 55370 2916
rect 55493 2907 55551 2913
rect 55493 2873 55505 2907
rect 55539 2904 55551 2907
rect 56594 2904 56600 2916
rect 55539 2876 56600 2904
rect 55539 2873 55551 2876
rect 55493 2867 55551 2873
rect 56594 2864 56600 2876
rect 56652 2864 56658 2916
rect 58526 2864 58532 2916
rect 58584 2864 58590 2916
rect 62117 2907 62175 2913
rect 62117 2873 62129 2907
rect 62163 2904 62175 2907
rect 62574 2904 62580 2916
rect 62163 2876 62580 2904
rect 62163 2873 62175 2876
rect 62117 2867 62175 2873
rect 62574 2864 62580 2876
rect 62632 2864 62638 2916
rect 47452 2808 49648 2836
rect 47452 2796 47458 2808
rect 51074 2796 51080 2848
rect 51132 2796 51138 2848
rect 51166 2796 51172 2848
rect 51224 2796 51230 2848
rect 54757 2839 54815 2845
rect 54757 2805 54769 2839
rect 54803 2836 54815 2839
rect 55214 2836 55220 2848
rect 54803 2808 55220 2836
rect 54803 2805 54815 2808
rect 54757 2799 54815 2805
rect 55214 2796 55220 2808
rect 55272 2796 55278 2848
rect 56229 2839 56287 2845
rect 56229 2805 56241 2839
rect 56275 2836 56287 2839
rect 56870 2836 56876 2848
rect 56275 2808 56876 2836
rect 56275 2805 56287 2808
rect 56229 2799 56287 2805
rect 56870 2796 56876 2808
rect 56928 2796 56934 2848
rect 56962 2796 56968 2848
rect 57020 2796 57026 2848
rect 58437 2839 58495 2845
rect 58437 2805 58449 2839
rect 58483 2836 58495 2839
rect 58894 2836 58900 2848
rect 58483 2808 58900 2836
rect 58483 2805 58495 2808
rect 58437 2799 58495 2805
rect 58894 2796 58900 2808
rect 58952 2796 58958 2848
rect 59906 2796 59912 2848
rect 59964 2796 59970 2848
rect 60645 2839 60703 2845
rect 60645 2805 60657 2839
rect 60691 2836 60703 2839
rect 61102 2836 61108 2848
rect 60691 2808 61108 2836
rect 60691 2805 60703 2808
rect 60645 2799 60703 2805
rect 61102 2796 61108 2808
rect 61160 2796 61166 2848
rect 64601 2839 64659 2845
rect 64601 2805 64613 2839
rect 64647 2836 64659 2839
rect 64966 2836 64972 2848
rect 64647 2808 64972 2836
rect 64647 2805 64659 2808
rect 64601 2799 64659 2805
rect 64966 2796 64972 2808
rect 65024 2796 65030 2848
rect 65720 2836 65748 2935
rect 67192 2904 67220 2935
rect 69014 2932 69020 2984
rect 69072 2932 69078 2984
rect 69474 2932 69480 2984
rect 69532 2972 69538 2984
rect 69661 2975 69719 2981
rect 69661 2972 69673 2975
rect 69532 2944 69673 2972
rect 69532 2932 69538 2944
rect 69661 2941 69673 2944
rect 69707 2941 69719 2975
rect 69661 2935 69719 2941
rect 71038 2932 71044 2984
rect 71096 2932 71102 2984
rect 71317 2975 71375 2981
rect 71317 2941 71329 2975
rect 71363 2972 71375 2975
rect 73246 2972 73252 2984
rect 71363 2944 73252 2972
rect 71363 2941 71375 2944
rect 71317 2935 71375 2941
rect 73246 2932 73252 2944
rect 73304 2932 73310 2984
rect 69382 2904 69388 2916
rect 67192 2876 69388 2904
rect 69382 2864 69388 2876
rect 69440 2864 69446 2916
rect 70305 2907 70363 2913
rect 70305 2873 70317 2907
rect 70351 2904 70363 2907
rect 70670 2904 70676 2916
rect 70351 2876 70676 2904
rect 70351 2873 70363 2876
rect 70305 2867 70363 2873
rect 70670 2864 70676 2876
rect 70728 2864 70734 2916
rect 66254 2836 66260 2848
rect 65720 2808 66260 2836
rect 66254 2796 66260 2808
rect 66312 2796 66318 2848
rect 66990 2796 66996 2848
rect 67048 2796 67054 2848
rect 67729 2839 67787 2845
rect 67729 2805 67741 2839
rect 67775 2836 67787 2839
rect 68462 2836 68468 2848
rect 67775 2808 68468 2836
rect 67775 2805 67787 2808
rect 67729 2799 67787 2805
rect 68462 2796 68468 2808
rect 68520 2796 68526 2848
rect 70397 2839 70455 2845
rect 70397 2805 70409 2839
rect 70443 2836 70455 2839
rect 70854 2836 70860 2848
rect 70443 2808 70860 2836
rect 70443 2805 70455 2808
rect 70397 2799 70455 2805
rect 70854 2796 70860 2808
rect 70912 2796 70918 2848
rect 71869 2839 71927 2845
rect 71869 2805 71881 2839
rect 71915 2836 71927 2839
rect 72234 2836 72240 2848
rect 71915 2808 72240 2836
rect 71915 2805 71927 2808
rect 71869 2799 71927 2805
rect 72234 2796 72240 2808
rect 72292 2796 72298 2848
rect 1012 2746 74980 2768
rect 1012 2694 1858 2746
rect 1910 2694 1922 2746
rect 1974 2694 1986 2746
rect 2038 2694 2050 2746
rect 2102 2694 2114 2746
rect 2166 2694 11858 2746
rect 11910 2694 11922 2746
rect 11974 2694 11986 2746
rect 12038 2694 12050 2746
rect 12102 2694 12114 2746
rect 12166 2694 21858 2746
rect 21910 2694 21922 2746
rect 21974 2694 21986 2746
rect 22038 2694 22050 2746
rect 22102 2694 22114 2746
rect 22166 2694 31858 2746
rect 31910 2694 31922 2746
rect 31974 2694 31986 2746
rect 32038 2694 32050 2746
rect 32102 2694 32114 2746
rect 32166 2694 41858 2746
rect 41910 2694 41922 2746
rect 41974 2694 41986 2746
rect 42038 2694 42050 2746
rect 42102 2694 42114 2746
rect 42166 2694 51858 2746
rect 51910 2694 51922 2746
rect 51974 2694 51986 2746
rect 52038 2694 52050 2746
rect 52102 2694 52114 2746
rect 52166 2694 61858 2746
rect 61910 2694 61922 2746
rect 61974 2694 61986 2746
rect 62038 2694 62050 2746
rect 62102 2694 62114 2746
rect 62166 2694 71858 2746
rect 71910 2694 71922 2746
rect 71974 2694 71986 2746
rect 72038 2694 72050 2746
rect 72102 2694 72114 2746
rect 72166 2694 74980 2746
rect 1012 2672 74980 2694
rect 22649 2635 22707 2641
rect 22649 2601 22661 2635
rect 22695 2632 22707 2635
rect 23106 2632 23112 2644
rect 22695 2604 23112 2632
rect 22695 2601 22707 2604
rect 22649 2595 22707 2601
rect 23106 2592 23112 2604
rect 23164 2592 23170 2644
rect 23385 2635 23443 2641
rect 23385 2601 23397 2635
rect 23431 2632 23443 2635
rect 23842 2632 23848 2644
rect 23431 2604 23848 2632
rect 23431 2601 23443 2604
rect 23385 2595 23443 2601
rect 23842 2592 23848 2604
rect 23900 2592 23906 2644
rect 26697 2635 26755 2641
rect 23952 2604 24532 2632
rect 22833 2499 22891 2505
rect 22833 2465 22845 2499
rect 22879 2496 22891 2499
rect 23952 2496 23980 2604
rect 24026 2524 24032 2576
rect 24084 2524 24090 2576
rect 22879 2468 23980 2496
rect 24044 2496 24072 2524
rect 24044 2468 24348 2496
rect 22879 2465 22891 2468
rect 22833 2459 22891 2465
rect 22097 2431 22155 2437
rect 22097 2397 22109 2431
rect 22143 2428 22155 2431
rect 24026 2428 24032 2440
rect 22143 2400 24032 2428
rect 22143 2397 22155 2400
rect 22097 2391 22155 2397
rect 24026 2388 24032 2400
rect 24084 2388 24090 2440
rect 24320 2437 24348 2468
rect 24121 2431 24179 2437
rect 24121 2397 24133 2431
rect 24167 2397 24179 2431
rect 24121 2391 24179 2397
rect 24305 2431 24363 2437
rect 24305 2397 24317 2431
rect 24351 2397 24363 2431
rect 24504 2428 24532 2604
rect 26697 2601 26709 2635
rect 26743 2632 26755 2635
rect 27706 2632 27712 2644
rect 26743 2604 27712 2632
rect 26743 2601 26755 2604
rect 26697 2595 26755 2601
rect 27706 2592 27712 2604
rect 27764 2592 27770 2644
rect 27982 2592 27988 2644
rect 28040 2632 28046 2644
rect 28261 2635 28319 2641
rect 28261 2632 28273 2635
rect 28040 2604 28273 2632
rect 28040 2592 28046 2604
rect 28261 2601 28273 2604
rect 28307 2601 28319 2635
rect 28261 2595 28319 2601
rect 29362 2592 29368 2644
rect 29420 2632 29426 2644
rect 29457 2635 29515 2641
rect 29457 2632 29469 2635
rect 29420 2604 29469 2632
rect 29420 2592 29426 2604
rect 29457 2601 29469 2604
rect 29503 2601 29515 2635
rect 29457 2595 29515 2601
rect 29546 2592 29552 2644
rect 29604 2632 29610 2644
rect 29641 2635 29699 2641
rect 29641 2632 29653 2635
rect 29604 2604 29653 2632
rect 29604 2592 29610 2604
rect 29641 2601 29653 2604
rect 29687 2601 29699 2635
rect 29641 2595 29699 2601
rect 30101 2635 30159 2641
rect 30101 2601 30113 2635
rect 30147 2632 30159 2635
rect 30466 2632 30472 2644
rect 30147 2604 30472 2632
rect 30147 2601 30159 2604
rect 30101 2595 30159 2601
rect 30466 2592 30472 2604
rect 30524 2592 30530 2644
rect 32217 2635 32275 2641
rect 32217 2601 32229 2635
rect 32263 2632 32275 2635
rect 32306 2632 32312 2644
rect 32263 2604 32312 2632
rect 32263 2601 32275 2604
rect 32217 2595 32275 2601
rect 32306 2592 32312 2604
rect 32364 2592 32370 2644
rect 34425 2635 34483 2641
rect 34425 2601 34437 2635
rect 34471 2632 34483 2635
rect 34606 2632 34612 2644
rect 34471 2604 34612 2632
rect 34471 2601 34483 2604
rect 34425 2595 34483 2601
rect 34606 2592 34612 2604
rect 34664 2592 34670 2644
rect 35437 2635 35495 2641
rect 35437 2601 35449 2635
rect 35483 2632 35495 2635
rect 36078 2632 36084 2644
rect 35483 2604 36084 2632
rect 35483 2601 35495 2604
rect 35437 2595 35495 2601
rect 36078 2592 36084 2604
rect 36136 2592 36142 2644
rect 36906 2592 36912 2644
rect 36964 2592 36970 2644
rect 37645 2635 37703 2641
rect 37645 2601 37657 2635
rect 37691 2632 37703 2635
rect 38378 2632 38384 2644
rect 37691 2604 38384 2632
rect 37691 2601 37703 2604
rect 37645 2595 37703 2601
rect 38378 2592 38384 2604
rect 38436 2592 38442 2644
rect 40218 2592 40224 2644
rect 40276 2632 40282 2644
rect 41233 2635 41291 2641
rect 41233 2632 41245 2635
rect 40276 2604 41245 2632
rect 40276 2592 40282 2604
rect 41233 2601 41245 2604
rect 41279 2601 41291 2635
rect 41233 2595 41291 2601
rect 42978 2592 42984 2644
rect 43036 2632 43042 2644
rect 43349 2635 43407 2641
rect 43349 2632 43361 2635
rect 43036 2604 43361 2632
rect 43036 2592 43042 2604
rect 43349 2601 43361 2604
rect 43395 2601 43407 2635
rect 43349 2595 43407 2601
rect 44634 2592 44640 2644
rect 44692 2632 44698 2644
rect 44913 2635 44971 2641
rect 44913 2632 44925 2635
rect 44692 2604 44925 2632
rect 44692 2592 44698 2604
rect 44913 2601 44925 2604
rect 44959 2601 44971 2635
rect 44913 2595 44971 2601
rect 45554 2592 45560 2644
rect 45612 2632 45618 2644
rect 45649 2635 45707 2641
rect 45649 2632 45661 2635
rect 45612 2604 45661 2632
rect 45612 2592 45618 2604
rect 45649 2601 45661 2604
rect 45695 2601 45707 2635
rect 45649 2595 45707 2601
rect 46106 2592 46112 2644
rect 46164 2632 46170 2644
rect 46385 2635 46443 2641
rect 46385 2632 46397 2635
rect 46164 2604 46397 2632
rect 46164 2592 46170 2604
rect 46385 2601 46397 2604
rect 46431 2601 46443 2635
rect 46385 2595 46443 2601
rect 48593 2635 48651 2641
rect 48593 2601 48605 2635
rect 48639 2632 48651 2635
rect 48774 2632 48780 2644
rect 48639 2604 48780 2632
rect 48639 2601 48651 2604
rect 48593 2595 48651 2601
rect 48774 2592 48780 2604
rect 48832 2592 48838 2644
rect 49421 2635 49479 2641
rect 49421 2601 49433 2635
rect 49467 2632 49479 2635
rect 49510 2632 49516 2644
rect 49467 2604 49516 2632
rect 49467 2601 49479 2604
rect 49421 2595 49479 2601
rect 49510 2592 49516 2604
rect 49568 2592 49574 2644
rect 50706 2592 50712 2644
rect 50764 2632 50770 2644
rect 50801 2635 50859 2641
rect 50801 2632 50813 2635
rect 50764 2604 50813 2632
rect 50764 2592 50770 2604
rect 50801 2601 50813 2604
rect 50847 2601 50859 2635
rect 50801 2595 50859 2601
rect 51534 2592 51540 2644
rect 51592 2592 51598 2644
rect 53006 2592 53012 2644
rect 53064 2592 53070 2644
rect 54757 2635 54815 2641
rect 54757 2601 54769 2635
rect 54803 2632 54815 2635
rect 54803 2604 64874 2632
rect 54803 2601 54815 2604
rect 54757 2595 54815 2601
rect 26602 2564 26608 2576
rect 24688 2536 26608 2564
rect 24688 2505 24716 2536
rect 26602 2524 26608 2536
rect 26660 2524 26666 2576
rect 30006 2524 30012 2576
rect 30064 2524 30070 2576
rect 31481 2567 31539 2573
rect 31481 2533 31493 2567
rect 31527 2564 31539 2567
rect 32674 2564 32680 2576
rect 31527 2536 32680 2564
rect 31527 2533 31539 2536
rect 31481 2527 31539 2533
rect 32674 2524 32680 2536
rect 32732 2524 32738 2576
rect 33689 2567 33747 2573
rect 33689 2533 33701 2567
rect 33735 2564 33747 2567
rect 34698 2564 34704 2576
rect 33735 2536 34704 2564
rect 33735 2533 33747 2536
rect 33689 2527 33747 2533
rect 34698 2524 34704 2536
rect 34756 2524 34762 2576
rect 34790 2524 34796 2576
rect 34848 2564 34854 2576
rect 54662 2564 54668 2576
rect 34848 2536 54668 2564
rect 34848 2524 34854 2536
rect 54662 2524 54668 2536
rect 54720 2524 54726 2576
rect 55950 2524 55956 2576
rect 56008 2524 56014 2576
rect 59817 2567 59875 2573
rect 59817 2533 59829 2567
rect 59863 2564 59875 2567
rect 60642 2564 60648 2576
rect 59863 2536 60648 2564
rect 59863 2533 59875 2536
rect 59817 2527 59875 2533
rect 60642 2524 60648 2536
rect 60700 2524 60706 2576
rect 61562 2524 61568 2576
rect 61620 2564 61626 2576
rect 61841 2567 61899 2573
rect 61841 2564 61853 2567
rect 61620 2536 61853 2564
rect 61620 2524 61626 2536
rect 61841 2533 61853 2536
rect 61887 2533 61899 2567
rect 61841 2527 61899 2533
rect 63310 2524 63316 2576
rect 63368 2524 63374 2576
rect 64417 2567 64475 2573
rect 64417 2533 64429 2567
rect 64463 2564 64475 2567
rect 64690 2564 64696 2576
rect 64463 2536 64696 2564
rect 64463 2533 64475 2536
rect 64417 2527 64475 2533
rect 64690 2524 64696 2536
rect 64748 2524 64754 2576
rect 64846 2564 64874 2604
rect 65242 2592 65248 2644
rect 65300 2632 65306 2644
rect 65521 2635 65579 2641
rect 65521 2632 65533 2635
rect 65300 2604 65533 2632
rect 65300 2592 65306 2604
rect 65521 2601 65533 2604
rect 65567 2601 65579 2635
rect 65521 2595 65579 2601
rect 66254 2592 66260 2644
rect 66312 2592 66318 2644
rect 69106 2592 69112 2644
rect 69164 2592 69170 2644
rect 71038 2592 71044 2644
rect 71096 2632 71102 2644
rect 71409 2635 71467 2641
rect 71409 2632 71421 2635
rect 71096 2604 71421 2632
rect 71096 2592 71102 2604
rect 71409 2601 71421 2604
rect 71455 2601 71467 2635
rect 71409 2595 71467 2601
rect 69658 2564 69664 2576
rect 64846 2536 69664 2564
rect 69658 2524 69664 2536
rect 69716 2524 69722 2576
rect 71222 2564 71228 2576
rect 69768 2536 71228 2564
rect 24673 2499 24731 2505
rect 24673 2465 24685 2499
rect 24719 2465 24731 2499
rect 24673 2459 24731 2465
rect 25225 2499 25283 2505
rect 25225 2465 25237 2499
rect 25271 2496 25283 2499
rect 26053 2499 26111 2505
rect 26053 2496 26065 2499
rect 25271 2468 26065 2496
rect 25271 2465 25283 2468
rect 25225 2459 25283 2465
rect 26053 2465 26065 2468
rect 26099 2465 26111 2499
rect 26053 2459 26111 2465
rect 28721 2499 28779 2505
rect 28721 2465 28733 2499
rect 28767 2496 28779 2499
rect 30098 2496 30104 2508
rect 28767 2468 30104 2496
rect 28767 2465 28779 2468
rect 28721 2459 28779 2465
rect 30098 2456 30104 2468
rect 30156 2456 30162 2508
rect 30742 2456 30748 2508
rect 30800 2456 30806 2508
rect 30929 2499 30987 2505
rect 30929 2465 30941 2499
rect 30975 2496 30987 2499
rect 31110 2496 31116 2508
rect 30975 2468 31116 2496
rect 30975 2465 30987 2468
rect 30929 2459 30987 2465
rect 31110 2456 31116 2468
rect 31168 2456 31174 2508
rect 31665 2499 31723 2505
rect 31665 2465 31677 2499
rect 31711 2496 31723 2499
rect 32398 2496 32404 2508
rect 31711 2468 32404 2496
rect 31711 2465 31723 2468
rect 31665 2459 31723 2465
rect 32398 2456 32404 2468
rect 32456 2456 32462 2508
rect 33778 2456 33784 2508
rect 33836 2456 33842 2508
rect 34885 2499 34943 2505
rect 34885 2465 34897 2499
rect 34931 2496 34943 2499
rect 34931 2468 35894 2496
rect 34931 2465 34943 2468
rect 34885 2459 34943 2465
rect 24504 2400 25360 2428
rect 24305 2391 24363 2397
rect 24136 2360 24164 2391
rect 24578 2360 24584 2372
rect 24136 2332 24584 2360
rect 24578 2320 24584 2332
rect 24636 2320 24642 2372
rect 25332 2360 25360 2400
rect 25406 2388 25412 2440
rect 25464 2388 25470 2440
rect 27062 2428 27068 2440
rect 26206 2400 27068 2428
rect 26206 2360 26234 2400
rect 27062 2388 27068 2400
rect 27120 2388 27126 2440
rect 28169 2431 28227 2437
rect 28169 2397 28181 2431
rect 28215 2428 28227 2431
rect 28258 2428 28264 2440
rect 28215 2400 28264 2428
rect 28215 2397 28227 2400
rect 28169 2391 28227 2397
rect 28258 2388 28264 2400
rect 28316 2388 28322 2440
rect 28442 2388 28448 2440
rect 28500 2388 28506 2440
rect 29273 2431 29331 2437
rect 29273 2397 29285 2431
rect 29319 2428 29331 2431
rect 31018 2428 31024 2440
rect 29319 2400 31024 2428
rect 29319 2397 29331 2400
rect 29273 2391 29331 2397
rect 31018 2388 31024 2400
rect 31076 2388 31082 2440
rect 32309 2431 32367 2437
rect 32309 2397 32321 2431
rect 32355 2397 32367 2431
rect 32309 2391 32367 2397
rect 25332 2332 26234 2360
rect 26786 2320 26792 2372
rect 26844 2360 26850 2372
rect 26973 2363 27031 2369
rect 26973 2360 26985 2363
rect 26844 2332 26985 2360
rect 26844 2320 26850 2332
rect 26973 2329 26985 2332
rect 27019 2329 27031 2363
rect 26973 2323 27031 2329
rect 27522 2320 27528 2372
rect 27580 2360 27586 2372
rect 28902 2360 28908 2372
rect 27580 2332 28908 2360
rect 27580 2320 27586 2332
rect 28902 2320 28908 2332
rect 28960 2360 28966 2372
rect 29641 2363 29699 2369
rect 29641 2360 29653 2363
rect 28960 2332 29653 2360
rect 28960 2320 28966 2332
rect 29641 2329 29653 2332
rect 29687 2329 29699 2363
rect 32324 2360 32352 2391
rect 33042 2388 33048 2440
rect 33100 2388 33106 2440
rect 35526 2388 35532 2440
rect 35584 2388 35590 2440
rect 35866 2428 35894 2468
rect 36170 2456 36176 2508
rect 36228 2496 36234 2508
rect 36265 2499 36323 2505
rect 36265 2496 36277 2499
rect 36228 2468 36277 2496
rect 36228 2456 36234 2468
rect 36265 2465 36277 2468
rect 36311 2465 36323 2499
rect 36265 2459 36323 2465
rect 37826 2456 37832 2508
rect 37884 2496 37890 2508
rect 38381 2499 38439 2505
rect 38381 2496 38393 2499
rect 37884 2468 38393 2496
rect 37884 2456 37890 2468
rect 38381 2465 38393 2468
rect 38427 2465 38439 2499
rect 38381 2459 38439 2465
rect 38746 2456 38752 2508
rect 38804 2456 38810 2508
rect 41506 2456 41512 2508
rect 41564 2496 41570 2508
rect 41785 2499 41843 2505
rect 41785 2496 41797 2499
rect 41564 2468 41797 2496
rect 41564 2456 41570 2468
rect 41785 2465 41797 2468
rect 41831 2465 41843 2499
rect 41785 2459 41843 2465
rect 42518 2456 42524 2508
rect 42576 2496 42582 2508
rect 42705 2499 42763 2505
rect 42705 2496 42717 2499
rect 42576 2468 42717 2496
rect 42576 2456 42582 2468
rect 42705 2465 42717 2468
rect 42751 2465 42763 2499
rect 42705 2459 42763 2465
rect 43438 2456 43444 2508
rect 43496 2456 43502 2508
rect 46934 2456 46940 2508
rect 46992 2456 46998 2508
rect 47118 2456 47124 2508
rect 47176 2456 47182 2508
rect 47302 2456 47308 2508
rect 47360 2496 47366 2508
rect 49786 2496 49792 2508
rect 47360 2468 49792 2496
rect 47360 2456 47366 2468
rect 49786 2456 49792 2468
rect 49844 2456 49850 2508
rect 49970 2456 49976 2508
rect 50028 2496 50034 2508
rect 50617 2499 50675 2505
rect 50617 2496 50629 2499
rect 50028 2468 50629 2496
rect 50028 2456 50034 2468
rect 50617 2465 50629 2468
rect 50663 2465 50675 2499
rect 50617 2459 50675 2465
rect 51074 2456 51080 2508
rect 51132 2496 51138 2508
rect 52089 2499 52147 2505
rect 52089 2496 52101 2499
rect 51132 2468 52101 2496
rect 51132 2456 51138 2468
rect 52089 2465 52101 2468
rect 52135 2465 52147 2499
rect 52089 2459 52147 2465
rect 54018 2456 54024 2508
rect 54076 2496 54082 2508
rect 54297 2499 54355 2505
rect 54297 2496 54309 2499
rect 54076 2468 54309 2496
rect 54076 2456 54082 2468
rect 54297 2465 54309 2468
rect 54343 2465 54355 2499
rect 54297 2459 54355 2465
rect 55214 2456 55220 2508
rect 55272 2456 55278 2508
rect 56594 2456 56600 2508
rect 56652 2456 56658 2508
rect 56870 2456 56876 2508
rect 56928 2496 56934 2508
rect 57241 2499 57299 2505
rect 57241 2496 57253 2499
rect 56928 2468 57253 2496
rect 56928 2456 56934 2468
rect 57241 2465 57253 2468
rect 57287 2465 57299 2499
rect 57241 2459 57299 2465
rect 58894 2456 58900 2508
rect 58952 2456 58958 2508
rect 59906 2456 59912 2508
rect 59964 2496 59970 2508
rect 60369 2499 60427 2505
rect 60369 2496 60381 2499
rect 59964 2468 60381 2496
rect 59964 2456 59970 2468
rect 60369 2465 60381 2468
rect 60415 2465 60427 2499
rect 60369 2459 60427 2465
rect 61102 2456 61108 2508
rect 61160 2456 61166 2508
rect 61212 2468 62528 2496
rect 36354 2428 36360 2440
rect 35866 2400 36360 2428
rect 36354 2388 36360 2400
rect 36412 2388 36418 2440
rect 37093 2431 37151 2437
rect 37093 2397 37105 2431
rect 37139 2428 37151 2431
rect 37642 2428 37648 2440
rect 37139 2400 37648 2428
rect 37139 2397 37151 2400
rect 37093 2391 37151 2397
rect 37642 2388 37648 2400
rect 37700 2388 37706 2440
rect 37737 2431 37795 2437
rect 37737 2397 37749 2431
rect 37783 2397 37795 2431
rect 37737 2391 37795 2397
rect 40405 2431 40463 2437
rect 40405 2397 40417 2431
rect 40451 2428 40463 2431
rect 40497 2431 40555 2437
rect 40497 2428 40509 2431
rect 40451 2400 40509 2428
rect 40451 2397 40463 2400
rect 40405 2391 40463 2397
rect 40497 2397 40509 2400
rect 40543 2397 40555 2431
rect 40497 2391 40555 2397
rect 34606 2360 34612 2372
rect 32324 2332 34612 2360
rect 29641 2323 29699 2329
rect 34606 2320 34612 2332
rect 34664 2320 34670 2372
rect 36262 2320 36268 2372
rect 36320 2360 36326 2372
rect 37752 2360 37780 2391
rect 41046 2388 41052 2440
rect 41104 2388 41110 2440
rect 41969 2431 42027 2437
rect 41969 2397 41981 2431
rect 42015 2397 42027 2431
rect 41969 2391 42027 2397
rect 44085 2431 44143 2437
rect 44085 2397 44097 2431
rect 44131 2428 44143 2431
rect 44177 2431 44235 2437
rect 44177 2428 44189 2431
rect 44131 2400 44189 2428
rect 44131 2397 44143 2400
rect 44085 2391 44143 2397
rect 44177 2397 44189 2400
rect 44223 2397 44235 2431
rect 44177 2391 44235 2397
rect 36320 2332 37780 2360
rect 36320 2320 36326 2332
rect 40770 2320 40776 2372
rect 40828 2360 40834 2372
rect 41984 2360 42012 2391
rect 45554 2388 45560 2440
rect 45612 2388 45618 2440
rect 46106 2388 46112 2440
rect 46164 2428 46170 2440
rect 46201 2431 46259 2437
rect 46201 2428 46213 2431
rect 46164 2400 46213 2428
rect 46164 2388 46170 2400
rect 46201 2397 46213 2400
rect 46247 2397 46259 2431
rect 46201 2391 46259 2397
rect 47765 2431 47823 2437
rect 47765 2397 47777 2431
rect 47811 2428 47823 2431
rect 47857 2431 47915 2437
rect 47857 2428 47869 2431
rect 47811 2400 47869 2428
rect 47811 2397 47823 2400
rect 47765 2391 47823 2397
rect 47857 2397 47869 2400
rect 47903 2397 47915 2431
rect 47857 2391 47915 2397
rect 49237 2431 49295 2437
rect 49237 2397 49249 2431
rect 49283 2428 49295 2431
rect 49418 2428 49424 2440
rect 49283 2400 49424 2428
rect 49283 2397 49295 2400
rect 49237 2391 49295 2397
rect 49418 2388 49424 2400
rect 49476 2388 49482 2440
rect 49605 2431 49663 2437
rect 49605 2397 49617 2431
rect 49651 2428 49663 2431
rect 50065 2431 50123 2437
rect 50065 2428 50077 2431
rect 49651 2400 50077 2428
rect 49651 2397 49663 2400
rect 49605 2391 49663 2397
rect 50065 2397 50077 2400
rect 50111 2397 50123 2431
rect 50065 2391 50123 2397
rect 51350 2388 51356 2440
rect 51408 2388 51414 2440
rect 51442 2388 51448 2440
rect 51500 2428 51506 2440
rect 52273 2431 52331 2437
rect 52273 2428 52285 2431
rect 51500 2400 52285 2428
rect 51500 2388 51506 2400
rect 52273 2397 52285 2400
rect 52319 2397 52331 2431
rect 52273 2391 52331 2397
rect 53653 2431 53711 2437
rect 53653 2397 53665 2431
rect 53699 2428 53711 2431
rect 53745 2431 53803 2437
rect 53745 2428 53757 2431
rect 53699 2400 53757 2428
rect 53699 2397 53711 2400
rect 53653 2391 53711 2397
rect 53745 2397 53757 2400
rect 53791 2397 53803 2431
rect 53745 2391 53803 2397
rect 54849 2431 54907 2437
rect 54849 2397 54861 2431
rect 54895 2428 54907 2431
rect 56686 2428 56692 2440
rect 54895 2400 56692 2428
rect 54895 2397 54907 2400
rect 54849 2391 54907 2397
rect 56686 2388 56692 2400
rect 56744 2388 56750 2440
rect 57517 2431 57575 2437
rect 57517 2397 57529 2431
rect 57563 2428 57575 2431
rect 58161 2431 58219 2437
rect 58161 2428 58173 2431
rect 57563 2400 58173 2428
rect 57563 2397 57575 2400
rect 57517 2391 57575 2397
rect 58161 2397 58173 2400
rect 58207 2397 58219 2431
rect 58161 2391 58219 2397
rect 58434 2388 58440 2440
rect 58492 2428 58498 2440
rect 58713 2431 58771 2437
rect 58713 2428 58725 2431
rect 58492 2400 58725 2428
rect 58492 2388 58498 2400
rect 58713 2397 58725 2400
rect 58759 2397 58771 2431
rect 58713 2391 58771 2397
rect 59722 2388 59728 2440
rect 59780 2428 59786 2440
rect 61212 2428 61240 2468
rect 59780 2400 61240 2428
rect 59780 2388 59786 2400
rect 61562 2388 61568 2440
rect 61620 2428 61626 2440
rect 62393 2431 62451 2437
rect 62393 2428 62405 2431
rect 61620 2400 62405 2428
rect 61620 2388 61626 2400
rect 62393 2397 62405 2400
rect 62439 2397 62451 2431
rect 62393 2391 62451 2397
rect 40828 2332 42012 2360
rect 44453 2363 44511 2369
rect 40828 2320 40834 2332
rect 44453 2329 44465 2363
rect 44499 2360 44511 2363
rect 47210 2360 47216 2372
rect 44499 2332 47216 2360
rect 44499 2329 44511 2332
rect 44453 2323 44511 2329
rect 47210 2320 47216 2332
rect 47268 2320 47274 2372
rect 47670 2320 47676 2372
rect 47728 2360 47734 2372
rect 50154 2360 50160 2372
rect 47728 2332 50160 2360
rect 47728 2320 47734 2332
rect 50154 2320 50160 2332
rect 50212 2320 50218 2372
rect 55861 2363 55919 2369
rect 55861 2329 55873 2363
rect 55907 2360 55919 2363
rect 57238 2360 57244 2372
rect 55907 2332 57244 2360
rect 55907 2329 55919 2332
rect 55861 2323 55919 2329
rect 57238 2320 57244 2332
rect 57296 2320 57302 2372
rect 60001 2363 60059 2369
rect 60001 2329 60013 2363
rect 60047 2360 60059 2363
rect 61654 2360 61660 2372
rect 60047 2332 61660 2360
rect 60047 2329 60059 2332
rect 60001 2323 60059 2329
rect 61654 2320 61660 2332
rect 61712 2320 61718 2372
rect 62500 2360 62528 2468
rect 62574 2456 62580 2508
rect 62632 2456 62638 2508
rect 62666 2456 62672 2508
rect 62724 2496 62730 2508
rect 62724 2468 64920 2496
rect 62724 2456 62730 2468
rect 62758 2388 62764 2440
rect 62816 2428 62822 2440
rect 63865 2431 63923 2437
rect 63865 2428 63877 2431
rect 62816 2400 63877 2428
rect 62816 2388 62822 2400
rect 63865 2397 63877 2400
rect 63911 2397 63923 2431
rect 63865 2391 63923 2397
rect 64782 2360 64788 2372
rect 62500 2332 64788 2360
rect 64782 2320 64788 2332
rect 64840 2320 64846 2372
rect 64892 2360 64920 2468
rect 64966 2456 64972 2508
rect 65024 2456 65030 2508
rect 66809 2499 66867 2505
rect 66809 2496 66821 2499
rect 65352 2468 66821 2496
rect 65352 2440 65380 2468
rect 66809 2465 66821 2468
rect 66855 2465 66867 2499
rect 66809 2459 66867 2465
rect 66990 2456 66996 2508
rect 67048 2456 67054 2508
rect 68462 2456 68468 2508
rect 68520 2456 68526 2508
rect 65334 2388 65340 2440
rect 65392 2388 65398 2440
rect 66070 2388 66076 2440
rect 66128 2388 66134 2440
rect 67082 2388 67088 2440
rect 67140 2428 67146 2440
rect 67729 2431 67787 2437
rect 67729 2428 67741 2431
rect 67140 2400 67741 2428
rect 67140 2388 67146 2400
rect 67729 2397 67741 2400
rect 67775 2397 67787 2431
rect 67729 2391 67787 2397
rect 68370 2388 68376 2440
rect 68428 2428 68434 2440
rect 69201 2431 69259 2437
rect 69201 2428 69213 2431
rect 68428 2400 69213 2428
rect 68428 2388 68434 2400
rect 69201 2397 69213 2400
rect 69247 2397 69259 2431
rect 69201 2391 69259 2397
rect 69768 2360 69796 2536
rect 71222 2524 71228 2536
rect 71280 2524 71286 2576
rect 70118 2456 70124 2508
rect 70176 2456 70182 2508
rect 70670 2456 70676 2508
rect 70728 2456 70734 2508
rect 72234 2456 72240 2508
rect 72292 2456 72298 2508
rect 70397 2431 70455 2437
rect 70397 2397 70409 2431
rect 70443 2397 70455 2431
rect 70397 2391 70455 2397
rect 71317 2431 71375 2437
rect 71317 2397 71329 2431
rect 71363 2428 71375 2431
rect 71961 2431 72019 2437
rect 71961 2428 71973 2431
rect 71363 2400 71973 2428
rect 71363 2397 71375 2400
rect 71317 2391 71375 2397
rect 71961 2397 71973 2400
rect 72007 2397 72019 2431
rect 71961 2391 72019 2397
rect 64892 2332 69796 2360
rect 70412 2360 70440 2391
rect 72234 2360 72240 2372
rect 70412 2332 72240 2360
rect 72234 2320 72240 2332
rect 72292 2320 72298 2372
rect 23474 2252 23480 2304
rect 23532 2252 23538 2304
rect 24489 2295 24547 2301
rect 24489 2261 24501 2295
rect 24535 2292 24547 2295
rect 25314 2292 25320 2304
rect 24535 2264 25320 2292
rect 24535 2261 24547 2264
rect 24489 2255 24547 2261
rect 25314 2252 25320 2264
rect 25372 2252 25378 2304
rect 25961 2295 26019 2301
rect 25961 2261 25973 2295
rect 26007 2292 26019 2295
rect 28626 2292 28632 2304
rect 26007 2264 28632 2292
rect 26007 2261 26019 2264
rect 25961 2255 26019 2261
rect 28626 2252 28632 2264
rect 28684 2252 28690 2304
rect 32953 2295 33011 2301
rect 32953 2261 32965 2295
rect 32999 2292 33011 2295
rect 34882 2292 34888 2304
rect 32999 2264 34888 2292
rect 32999 2261 33011 2264
rect 32953 2255 33011 2261
rect 34882 2252 34888 2264
rect 34940 2252 34946 2304
rect 35710 2252 35716 2304
rect 35768 2292 35774 2304
rect 36173 2295 36231 2301
rect 36173 2292 36185 2295
rect 35768 2264 36185 2292
rect 35768 2252 35774 2264
rect 36173 2261 36185 2264
rect 36219 2261 36231 2295
rect 36173 2255 36231 2261
rect 39393 2295 39451 2301
rect 39393 2261 39405 2295
rect 39439 2292 39451 2295
rect 39574 2292 39580 2304
rect 39439 2264 39580 2292
rect 39439 2261 39451 2264
rect 39393 2255 39451 2261
rect 39574 2252 39580 2264
rect 39632 2252 39638 2304
rect 39761 2295 39819 2301
rect 39761 2261 39773 2295
rect 39807 2292 39819 2295
rect 40310 2292 40316 2304
rect 39807 2264 40316 2292
rect 39807 2261 39819 2264
rect 39761 2255 39819 2261
rect 40310 2252 40316 2264
rect 40368 2252 40374 2304
rect 42613 2295 42671 2301
rect 42613 2261 42625 2295
rect 42659 2292 42671 2295
rect 44818 2292 44824 2304
rect 42659 2264 44824 2292
rect 42659 2261 42671 2264
rect 42613 2255 42671 2261
rect 44818 2252 44824 2264
rect 44876 2252 44882 2304
rect 44910 2252 44916 2304
rect 44968 2292 44974 2304
rect 46934 2292 46940 2304
rect 44968 2264 46940 2292
rect 44968 2252 44974 2264
rect 46934 2252 46940 2264
rect 46992 2252 46998 2304
rect 48498 2252 48504 2304
rect 48556 2252 48562 2304
rect 52917 2295 52975 2301
rect 52917 2261 52929 2295
rect 52963 2292 52975 2295
rect 53190 2292 53196 2304
rect 52963 2264 53196 2292
rect 52963 2261 52975 2264
rect 52917 2255 52975 2261
rect 53190 2252 53196 2264
rect 53248 2252 53254 2304
rect 56042 2252 56048 2304
rect 56100 2292 56106 2304
rect 56689 2295 56747 2301
rect 56689 2292 56701 2295
rect 56100 2264 56701 2292
rect 56100 2252 56106 2264
rect 56689 2261 56701 2264
rect 56735 2261 56747 2295
rect 56689 2255 56747 2261
rect 58069 2295 58127 2301
rect 58069 2261 58081 2295
rect 58115 2292 58127 2295
rect 59446 2292 59452 2304
rect 58115 2264 59452 2292
rect 58115 2261 58127 2264
rect 58069 2255 58127 2261
rect 59446 2252 59452 2264
rect 59504 2252 59510 2304
rect 59538 2252 59544 2304
rect 59596 2252 59602 2304
rect 61013 2295 61071 2301
rect 61013 2261 61025 2295
rect 61059 2292 61071 2295
rect 61194 2292 61200 2304
rect 61059 2264 61200 2292
rect 61059 2261 61071 2264
rect 61013 2255 61071 2261
rect 61194 2252 61200 2264
rect 61252 2252 61258 2304
rect 61749 2295 61807 2301
rect 61749 2261 61761 2295
rect 61795 2292 61807 2295
rect 62482 2292 62488 2304
rect 61795 2264 62488 2292
rect 61795 2261 61807 2264
rect 61749 2255 61807 2261
rect 62482 2252 62488 2264
rect 62540 2252 62546 2304
rect 63221 2295 63279 2301
rect 63221 2261 63233 2295
rect 63267 2292 63279 2295
rect 64966 2292 64972 2304
rect 63267 2264 64972 2292
rect 63267 2261 63279 2264
rect 63221 2255 63279 2261
rect 64966 2252 64972 2264
rect 65024 2252 65030 2304
rect 67637 2295 67695 2301
rect 67637 2261 67649 2295
rect 67683 2292 67695 2295
rect 68094 2292 68100 2304
rect 67683 2264 68100 2292
rect 67683 2261 67695 2264
rect 67637 2255 67695 2261
rect 68094 2252 68100 2264
rect 68152 2252 68158 2304
rect 68373 2295 68431 2301
rect 68373 2261 68385 2295
rect 68419 2292 68431 2295
rect 69750 2292 69756 2304
rect 68419 2264 69756 2292
rect 68419 2261 68431 2264
rect 68373 2255 68431 2261
rect 69750 2252 69756 2264
rect 69808 2252 69814 2304
rect 69845 2295 69903 2301
rect 69845 2261 69857 2295
rect 69891 2292 69903 2295
rect 70670 2292 70676 2304
rect 69891 2264 70676 2292
rect 69891 2261 69903 2264
rect 69845 2255 69903 2261
rect 70670 2252 70676 2264
rect 70728 2252 70734 2304
rect 72789 2295 72847 2301
rect 72789 2261 72801 2295
rect 72835 2292 72847 2295
rect 74626 2292 74632 2304
rect 72835 2264 74632 2292
rect 72835 2261 72847 2264
rect 72789 2255 72847 2261
rect 74626 2252 74632 2264
rect 74684 2252 74690 2304
rect 1012 2202 74980 2224
rect 1012 2150 4210 2202
rect 4262 2150 4274 2202
rect 4326 2150 4338 2202
rect 4390 2150 4402 2202
rect 4454 2150 4466 2202
rect 4518 2150 14210 2202
rect 14262 2150 14274 2202
rect 14326 2150 14338 2202
rect 14390 2150 14402 2202
rect 14454 2150 14466 2202
rect 14518 2150 24210 2202
rect 24262 2150 24274 2202
rect 24326 2150 24338 2202
rect 24390 2150 24402 2202
rect 24454 2150 24466 2202
rect 24518 2150 34210 2202
rect 34262 2150 34274 2202
rect 34326 2150 34338 2202
rect 34390 2150 34402 2202
rect 34454 2150 34466 2202
rect 34518 2150 44210 2202
rect 44262 2150 44274 2202
rect 44326 2150 44338 2202
rect 44390 2150 44402 2202
rect 44454 2150 44466 2202
rect 44518 2150 54210 2202
rect 54262 2150 54274 2202
rect 54326 2150 54338 2202
rect 54390 2150 54402 2202
rect 54454 2150 54466 2202
rect 54518 2150 64210 2202
rect 64262 2150 64274 2202
rect 64326 2150 64338 2202
rect 64390 2150 64402 2202
rect 64454 2150 64466 2202
rect 64518 2150 74210 2202
rect 74262 2150 74274 2202
rect 74326 2150 74338 2202
rect 74390 2150 74402 2202
rect 74454 2150 74466 2202
rect 74518 2150 74980 2202
rect 1012 2128 74980 2150
rect 21545 2091 21603 2097
rect 21545 2057 21557 2091
rect 21591 2088 21603 2091
rect 22370 2088 22376 2100
rect 21591 2060 22376 2088
rect 21591 2057 21603 2060
rect 21545 2051 21603 2057
rect 22370 2048 22376 2060
rect 22428 2048 22434 2100
rect 24946 2088 24952 2100
rect 22664 2060 24952 2088
rect 22189 1955 22247 1961
rect 22189 1921 22201 1955
rect 22235 1952 22247 1955
rect 22664 1952 22692 2060
rect 24946 2048 24952 2060
rect 25004 2048 25010 2100
rect 25961 2091 26019 2097
rect 25961 2057 25973 2091
rect 26007 2088 26019 2091
rect 26234 2088 26240 2100
rect 26007 2060 26240 2088
rect 26007 2057 26019 2060
rect 25961 2051 26019 2057
rect 26234 2048 26240 2060
rect 26292 2048 26298 2100
rect 26973 2091 27031 2097
rect 26973 2057 26985 2091
rect 27019 2088 27031 2091
rect 27614 2088 27620 2100
rect 27019 2060 27620 2088
rect 27019 2057 27031 2060
rect 26973 2051 27031 2057
rect 27614 2048 27620 2060
rect 27672 2048 27678 2100
rect 33318 2088 33324 2100
rect 30208 2060 33324 2088
rect 22741 2023 22799 2029
rect 22741 1989 22753 2023
rect 22787 2020 22799 2023
rect 22787 1992 24348 2020
rect 22787 1989 22799 1992
rect 22741 1983 22799 1989
rect 22235 1924 22692 1952
rect 22235 1921 22247 1924
rect 22189 1915 22247 1921
rect 23474 1912 23480 1964
rect 23532 1912 23538 1964
rect 24320 1961 24348 1992
rect 24305 1955 24363 1961
rect 24305 1921 24317 1955
rect 24351 1921 24363 1955
rect 24305 1915 24363 1921
rect 25222 1912 25228 1964
rect 25280 1952 25286 1964
rect 25777 1955 25835 1961
rect 25777 1952 25789 1955
rect 25280 1924 25789 1952
rect 25280 1912 25286 1924
rect 25777 1921 25789 1924
rect 25823 1921 25835 1955
rect 25777 1915 25835 1921
rect 26878 1912 26884 1964
rect 26936 1912 26942 1964
rect 26970 1912 26976 1964
rect 27028 1952 27034 1964
rect 27249 1955 27307 1961
rect 27249 1952 27261 1955
rect 27028 1924 27261 1952
rect 27028 1912 27034 1924
rect 27249 1921 27261 1924
rect 27295 1921 27307 1955
rect 27249 1915 27307 1921
rect 28994 1912 29000 1964
rect 29052 1912 29058 1964
rect 30208 1961 30236 2060
rect 33318 2048 33324 2060
rect 33376 2048 33382 2100
rect 36262 2048 36268 2100
rect 36320 2048 36326 2100
rect 37001 2091 37059 2097
rect 37001 2057 37013 2091
rect 37047 2088 37059 2091
rect 37274 2088 37280 2100
rect 37047 2060 37280 2088
rect 37047 2057 37059 2060
rect 37001 2051 37059 2057
rect 37274 2048 37280 2060
rect 37332 2048 37338 2100
rect 39025 2091 39083 2097
rect 39025 2057 39037 2091
rect 39071 2088 39083 2091
rect 39114 2088 39120 2100
rect 39071 2060 39120 2088
rect 39071 2057 39083 2060
rect 39025 2051 39083 2057
rect 39114 2048 39120 2060
rect 39172 2048 39178 2100
rect 39761 2091 39819 2097
rect 39761 2057 39773 2091
rect 39807 2088 39819 2091
rect 39850 2088 39856 2100
rect 39807 2060 39856 2088
rect 39807 2057 39819 2060
rect 39761 2051 39819 2057
rect 39850 2048 39856 2060
rect 39908 2048 39914 2100
rect 40586 2048 40592 2100
rect 40644 2088 40650 2100
rect 41233 2091 41291 2097
rect 41233 2088 41245 2091
rect 40644 2060 41245 2088
rect 40644 2048 40650 2060
rect 41233 2057 41245 2060
rect 41279 2057 41291 2091
rect 41233 2051 41291 2057
rect 45370 2048 45376 2100
rect 45428 2048 45434 2100
rect 46106 2048 46112 2100
rect 46164 2048 46170 2100
rect 55858 2088 55864 2100
rect 46216 2060 55864 2088
rect 36538 2020 36544 2032
rect 30300 1992 36544 2020
rect 30193 1955 30251 1961
rect 30193 1921 30205 1955
rect 30239 1921 30251 1955
rect 30193 1915 30251 1921
rect 20993 1887 21051 1893
rect 20993 1853 21005 1887
rect 21039 1853 21051 1887
rect 20993 1847 21051 1853
rect 21008 1816 21036 1847
rect 23566 1844 23572 1896
rect 23624 1844 23630 1896
rect 24026 1844 24032 1896
rect 24084 1884 24090 1896
rect 25314 1884 25320 1896
rect 24084 1856 25320 1884
rect 24084 1844 24090 1856
rect 25314 1844 25320 1856
rect 25372 1844 25378 1896
rect 25501 1887 25559 1893
rect 25501 1853 25513 1887
rect 25547 1884 25559 1887
rect 25590 1884 25596 1896
rect 25547 1856 25596 1884
rect 25547 1853 25559 1856
rect 25501 1847 25559 1853
rect 25590 1844 25596 1856
rect 25648 1844 25654 1896
rect 26142 1844 26148 1896
rect 26200 1844 26206 1896
rect 28445 1887 28503 1893
rect 28445 1853 28457 1887
rect 28491 1884 28503 1887
rect 30300 1884 30328 1992
rect 36538 1980 36544 1992
rect 36596 1980 36602 2032
rect 46216 2020 46244 2060
rect 55858 2048 55864 2060
rect 55916 2048 55922 2100
rect 55953 2091 56011 2097
rect 55953 2057 55965 2091
rect 55999 2088 56011 2091
rect 56502 2088 56508 2100
rect 55999 2060 56508 2088
rect 55999 2057 56011 2060
rect 55953 2051 56011 2057
rect 56502 2048 56508 2060
rect 56560 2048 56566 2100
rect 58434 2048 58440 2100
rect 58492 2048 58498 2100
rect 60366 2048 60372 2100
rect 60424 2088 60430 2100
rect 60461 2091 60519 2097
rect 60461 2088 60473 2091
rect 60424 2060 60473 2088
rect 60424 2048 60430 2060
rect 60461 2057 60473 2060
rect 60507 2057 60519 2091
rect 60461 2051 60519 2057
rect 61378 2048 61384 2100
rect 61436 2088 61442 2100
rect 61933 2091 61991 2097
rect 61933 2088 61945 2091
rect 61436 2060 61945 2088
rect 61436 2048 61442 2060
rect 61933 2057 61945 2060
rect 61979 2057 61991 2091
rect 61933 2051 61991 2057
rect 66070 2048 66076 2100
rect 66128 2048 66134 2100
rect 69014 2048 69020 2100
rect 69072 2088 69078 2100
rect 70121 2091 70179 2097
rect 70121 2088 70133 2091
rect 69072 2060 70133 2088
rect 69072 2048 69078 2060
rect 70121 2057 70133 2060
rect 70167 2057 70179 2091
rect 72326 2088 72332 2100
rect 70121 2051 70179 2057
rect 70228 2060 72332 2088
rect 38580 1992 46244 2020
rect 46768 1992 48268 2020
rect 31849 1955 31907 1961
rect 31849 1921 31861 1955
rect 31895 1952 31907 1955
rect 32858 1952 32864 1964
rect 31895 1924 32864 1952
rect 31895 1921 31907 1924
rect 31849 1915 31907 1921
rect 32858 1912 32864 1924
rect 32916 1912 32922 1964
rect 33689 1955 33747 1961
rect 33689 1921 33701 1955
rect 33735 1952 33747 1955
rect 34790 1952 34796 1964
rect 33735 1924 34796 1952
rect 33735 1921 33747 1924
rect 33689 1915 33747 1921
rect 34790 1912 34796 1924
rect 34848 1912 34854 1964
rect 35529 1955 35587 1961
rect 35529 1921 35541 1955
rect 35575 1952 35587 1955
rect 35618 1952 35624 1964
rect 35575 1924 35624 1952
rect 35575 1921 35587 1924
rect 35529 1915 35587 1921
rect 35618 1912 35624 1924
rect 35676 1912 35682 1964
rect 35710 1912 35716 1964
rect 35768 1912 35774 1964
rect 36449 1955 36507 1961
rect 36449 1921 36461 1955
rect 36495 1952 36507 1955
rect 37458 1952 37464 1964
rect 36495 1924 37464 1952
rect 36495 1921 36507 1924
rect 36449 1915 36507 1921
rect 37458 1912 37464 1924
rect 37516 1912 37522 1964
rect 38580 1961 38608 1992
rect 38565 1955 38623 1961
rect 38565 1921 38577 1955
rect 38611 1921 38623 1955
rect 38565 1915 38623 1921
rect 39574 1912 39580 1964
rect 39632 1912 39638 1964
rect 40310 1912 40316 1964
rect 40368 1912 40374 1964
rect 41414 1912 41420 1964
rect 41472 1952 41478 1964
rect 41785 1955 41843 1961
rect 41785 1952 41797 1955
rect 41472 1924 41797 1952
rect 41472 1912 41478 1924
rect 41785 1921 41797 1924
rect 41831 1921 41843 1955
rect 41785 1915 41843 1921
rect 43809 1955 43867 1961
rect 43809 1921 43821 1955
rect 43855 1952 43867 1955
rect 44910 1952 44916 1964
rect 43855 1924 44916 1952
rect 43855 1921 43867 1924
rect 43809 1915 43867 1921
rect 44910 1912 44916 1924
rect 44968 1912 44974 1964
rect 45281 1955 45339 1961
rect 45281 1921 45293 1955
rect 45327 1921 45339 1955
rect 45281 1915 45339 1921
rect 28491 1856 30328 1884
rect 28491 1853 28503 1856
rect 28445 1847 28503 1853
rect 30374 1844 30380 1896
rect 30432 1884 30438 1896
rect 30653 1887 30711 1893
rect 30653 1884 30665 1887
rect 30432 1856 30665 1884
rect 30432 1844 30438 1856
rect 30653 1853 30665 1856
rect 30699 1853 30711 1887
rect 30653 1847 30711 1853
rect 32214 1844 32220 1896
rect 32272 1884 32278 1896
rect 32493 1887 32551 1893
rect 32493 1884 32505 1887
rect 32272 1856 32505 1884
rect 32272 1844 32278 1856
rect 32493 1853 32505 1856
rect 32539 1853 32551 1887
rect 32493 1847 32551 1853
rect 34054 1844 34060 1896
rect 34112 1884 34118 1896
rect 34333 1887 34391 1893
rect 34333 1884 34345 1887
rect 34112 1856 34345 1884
rect 34112 1844 34118 1856
rect 34333 1853 34345 1856
rect 34379 1853 34391 1887
rect 34333 1847 34391 1853
rect 36814 1844 36820 1896
rect 36872 1884 36878 1896
rect 37369 1887 37427 1893
rect 37369 1884 37381 1887
rect 36872 1856 37381 1884
rect 36872 1844 36878 1856
rect 37369 1853 37381 1856
rect 37415 1853 37427 1887
rect 37369 1847 37427 1853
rect 39114 1844 39120 1896
rect 39172 1884 39178 1896
rect 41049 1887 41107 1893
rect 41049 1884 41061 1887
rect 39172 1856 41061 1884
rect 39172 1844 39178 1856
rect 41049 1853 41061 1856
rect 41095 1853 41107 1887
rect 41049 1847 41107 1853
rect 42334 1844 42340 1896
rect 42392 1884 42398 1896
rect 42613 1887 42671 1893
rect 42613 1884 42625 1887
rect 42392 1856 42625 1884
rect 42392 1844 42398 1856
rect 42613 1853 42625 1856
rect 42659 1853 42671 1887
rect 42613 1847 42671 1853
rect 43714 1844 43720 1896
rect 43772 1884 43778 1896
rect 44177 1887 44235 1893
rect 44177 1884 44189 1887
rect 43772 1856 44189 1884
rect 43772 1844 43778 1856
rect 44177 1853 44189 1856
rect 44223 1853 44235 1887
rect 45296 1884 45324 1915
rect 45922 1912 45928 1964
rect 45980 1912 45986 1964
rect 46768 1952 46796 1992
rect 46032 1924 46796 1952
rect 46032 1884 46060 1924
rect 46842 1912 46848 1964
rect 46900 1912 46906 1964
rect 47026 1912 47032 1964
rect 47084 1952 47090 1964
rect 47489 1955 47547 1961
rect 47489 1952 47501 1955
rect 47084 1924 47501 1952
rect 47084 1912 47090 1924
rect 47489 1921 47501 1924
rect 47535 1921 47547 1955
rect 47489 1915 47547 1921
rect 45296 1856 46060 1884
rect 44177 1847 44235 1853
rect 46658 1844 46664 1896
rect 46716 1844 46722 1896
rect 47854 1844 47860 1896
rect 47912 1884 47918 1896
rect 48133 1887 48191 1893
rect 48133 1884 48145 1887
rect 47912 1856 48145 1884
rect 47912 1844 47918 1856
rect 48133 1853 48145 1856
rect 48179 1853 48191 1887
rect 48133 1847 48191 1853
rect 24213 1819 24271 1825
rect 21008 1788 24164 1816
rect 22830 1708 22836 1760
rect 22888 1708 22894 1760
rect 24136 1748 24164 1788
rect 24213 1785 24225 1819
rect 24259 1816 24271 1819
rect 27798 1816 27804 1828
rect 24259 1788 27804 1816
rect 24259 1785 24271 1788
rect 24213 1779 24271 1785
rect 27798 1776 27804 1788
rect 27856 1776 27862 1828
rect 28258 1776 28264 1828
rect 28316 1816 28322 1828
rect 48240 1816 48268 1992
rect 49418 1980 49424 2032
rect 49476 1980 49482 2032
rect 50525 2023 50583 2029
rect 50525 1989 50537 2023
rect 50571 2020 50583 2023
rect 51166 2020 51172 2032
rect 50571 1992 51172 2020
rect 50571 1989 50583 1992
rect 50525 1983 50583 1989
rect 51166 1980 51172 1992
rect 51224 1980 51230 2032
rect 52454 2020 52460 2032
rect 51644 1992 52460 2020
rect 49329 1955 49387 1961
rect 49329 1921 49341 1955
rect 49375 1952 49387 1955
rect 49602 1952 49608 1964
rect 49375 1924 49608 1952
rect 49375 1921 49387 1924
rect 49329 1915 49387 1921
rect 49602 1912 49608 1924
rect 49660 1912 49666 1964
rect 49878 1912 49884 1964
rect 49936 1952 49942 1964
rect 49973 1955 50031 1961
rect 49973 1952 49985 1955
rect 49936 1924 49985 1952
rect 49936 1912 49942 1924
rect 49973 1921 49985 1924
rect 50019 1921 50031 1955
rect 49973 1915 50031 1921
rect 50157 1955 50215 1961
rect 50157 1921 50169 1955
rect 50203 1952 50215 1955
rect 51644 1952 51672 1992
rect 52454 1980 52460 1992
rect 52512 1980 52518 2032
rect 52638 1980 52644 2032
rect 52696 1980 52702 2032
rect 52748 1992 68232 2020
rect 50203 1924 51672 1952
rect 52089 1955 52147 1961
rect 50203 1921 50215 1924
rect 50157 1915 50215 1921
rect 52089 1921 52101 1955
rect 52135 1952 52147 1955
rect 52270 1952 52276 1964
rect 52135 1924 52276 1952
rect 52135 1921 52147 1924
rect 52089 1915 52147 1921
rect 52270 1912 52276 1924
rect 52328 1912 52334 1964
rect 50614 1844 50620 1896
rect 50672 1884 50678 1896
rect 50893 1887 50951 1893
rect 50893 1884 50905 1887
rect 50672 1856 50905 1884
rect 50672 1844 50678 1856
rect 50893 1853 50905 1856
rect 50939 1853 50951 1887
rect 50893 1847 50951 1853
rect 52748 1816 52776 1992
rect 53190 1912 53196 1964
rect 53248 1912 53254 1964
rect 54849 1955 54907 1961
rect 54849 1921 54861 1955
rect 54895 1921 54907 1955
rect 54849 1915 54907 1921
rect 53374 1844 53380 1896
rect 53432 1884 53438 1896
rect 53653 1887 53711 1893
rect 53653 1884 53665 1887
rect 53432 1856 53665 1884
rect 53432 1844 53438 1856
rect 53653 1853 53665 1856
rect 53699 1853 53711 1887
rect 54864 1884 54892 1915
rect 54938 1912 54944 1964
rect 54996 1912 55002 1964
rect 55306 1912 55312 1964
rect 55364 1952 55370 1964
rect 55493 1955 55551 1961
rect 55493 1952 55505 1955
rect 55364 1924 55505 1952
rect 55364 1912 55370 1924
rect 55493 1921 55505 1924
rect 55539 1921 55551 1955
rect 55493 1915 55551 1921
rect 56042 1912 56048 1964
rect 56100 1912 56106 1964
rect 57606 1912 57612 1964
rect 57664 1912 57670 1964
rect 60369 1955 60427 1961
rect 60369 1921 60381 1955
rect 60415 1952 60427 1955
rect 60458 1952 60464 1964
rect 60415 1924 60464 1952
rect 60415 1921 60427 1924
rect 60369 1915 60427 1921
rect 60458 1912 60464 1924
rect 60516 1912 60522 1964
rect 61194 1912 61200 1964
rect 61252 1912 61258 1964
rect 62482 1912 62488 1964
rect 62540 1912 62546 1964
rect 63313 1955 63371 1961
rect 63313 1921 63325 1955
rect 63359 1952 63371 1955
rect 63359 1924 64184 1952
rect 63359 1921 63371 1924
rect 63313 1915 63371 1921
rect 54864 1856 56088 1884
rect 53653 1847 53711 1853
rect 28316 1788 47808 1816
rect 48240 1788 52776 1816
rect 56060 1816 56088 1856
rect 56134 1844 56140 1896
rect 56192 1884 56198 1896
rect 56413 1887 56471 1893
rect 56413 1884 56425 1887
rect 56192 1856 56425 1884
rect 56192 1844 56198 1856
rect 56413 1853 56425 1856
rect 56459 1853 56471 1887
rect 56413 1847 56471 1853
rect 56962 1844 56968 1896
rect 57020 1884 57026 1896
rect 57793 1887 57851 1893
rect 57793 1884 57805 1887
rect 57020 1856 57805 1884
rect 57020 1844 57026 1856
rect 57793 1853 57805 1856
rect 57839 1853 57851 1887
rect 57793 1847 57851 1853
rect 58894 1844 58900 1896
rect 58952 1884 58958 1896
rect 59173 1887 59231 1893
rect 59173 1884 59185 1887
rect 58952 1856 59185 1884
rect 58952 1844 58958 1856
rect 59173 1853 59185 1856
rect 59219 1853 59231 1887
rect 59173 1847 59231 1853
rect 59538 1844 59544 1896
rect 59596 1884 59602 1896
rect 61013 1887 61071 1893
rect 61013 1884 61025 1887
rect 59596 1856 61025 1884
rect 59596 1844 59602 1856
rect 61013 1853 61025 1856
rect 61059 1853 61071 1887
rect 62666 1884 62672 1896
rect 61013 1847 61071 1853
rect 61120 1856 62672 1884
rect 61120 1816 61148 1856
rect 62666 1844 62672 1856
rect 62724 1844 62730 1896
rect 63034 1844 63040 1896
rect 63092 1884 63098 1896
rect 63589 1887 63647 1893
rect 63589 1884 63601 1887
rect 63092 1856 63601 1884
rect 63092 1844 63098 1856
rect 63589 1853 63601 1856
rect 63635 1853 63647 1887
rect 64156 1884 64184 1924
rect 64598 1912 64604 1964
rect 64656 1912 64662 1964
rect 64708 1924 66760 1952
rect 64708 1884 64736 1924
rect 64156 1856 64736 1884
rect 63589 1847 63647 1853
rect 64782 1844 64788 1896
rect 64840 1884 64846 1896
rect 65061 1887 65119 1893
rect 65061 1884 65073 1887
rect 64840 1856 65073 1884
rect 64840 1844 64846 1856
rect 65061 1853 65073 1856
rect 65107 1853 65119 1887
rect 65061 1847 65119 1853
rect 66625 1887 66683 1893
rect 66625 1853 66637 1887
rect 66671 1853 66683 1887
rect 66625 1847 66683 1853
rect 56060 1788 61148 1816
rect 61841 1819 61899 1825
rect 28316 1776 28322 1788
rect 24854 1748 24860 1760
rect 24136 1720 24860 1748
rect 24854 1708 24860 1720
rect 24912 1708 24918 1760
rect 26697 1751 26755 1757
rect 26697 1717 26709 1751
rect 26743 1748 26755 1751
rect 31386 1748 31392 1760
rect 26743 1720 31392 1748
rect 26743 1717 26755 1720
rect 26697 1711 26755 1717
rect 31386 1708 31392 1720
rect 31444 1708 31450 1760
rect 40494 1708 40500 1760
rect 40552 1708 40558 1760
rect 43254 1708 43260 1760
rect 43312 1748 43318 1760
rect 46658 1748 46664 1760
rect 43312 1720 46664 1748
rect 43312 1708 43318 1720
rect 46658 1708 46664 1720
rect 46716 1708 46722 1760
rect 47029 1751 47087 1757
rect 47029 1717 47041 1751
rect 47075 1748 47087 1751
rect 47302 1748 47308 1760
rect 47075 1720 47308 1748
rect 47075 1717 47087 1720
rect 47029 1711 47087 1717
rect 47302 1708 47308 1720
rect 47360 1708 47366 1760
rect 47670 1708 47676 1760
rect 47728 1708 47734 1760
rect 47780 1748 47808 1788
rect 61841 1785 61853 1819
rect 61887 1816 61899 1819
rect 62390 1816 62396 1828
rect 61887 1788 62396 1816
rect 61887 1785 61899 1788
rect 61841 1779 61899 1785
rect 62390 1776 62396 1788
rect 62448 1776 62454 1828
rect 63954 1776 63960 1828
rect 64012 1816 64018 1828
rect 66640 1816 66668 1847
rect 64012 1788 66668 1816
rect 66732 1816 66760 1924
rect 66806 1912 66812 1964
rect 66864 1912 66870 1964
rect 68094 1912 68100 1964
rect 68152 1912 68158 1964
rect 68204 1952 68232 1992
rect 68278 1980 68284 2032
rect 68336 2020 68342 2032
rect 68373 2023 68431 2029
rect 68373 2020 68385 2023
rect 68336 1992 68385 2020
rect 68336 1980 68342 1992
rect 68373 1989 68385 1992
rect 68419 1989 68431 2023
rect 70228 2020 70256 2060
rect 72326 2048 72332 2060
rect 72384 2048 72390 2100
rect 68373 1983 68431 1989
rect 68480 1992 70256 2020
rect 68480 1952 68508 1992
rect 71130 1980 71136 2032
rect 71188 1980 71194 2032
rect 73430 1980 73436 2032
rect 73488 1980 73494 2032
rect 68204 1924 68508 1952
rect 68646 1912 68652 1964
rect 68704 1912 68710 1964
rect 70670 1912 70676 1964
rect 70728 1912 70734 1964
rect 70854 1912 70860 1964
rect 70912 1912 70918 1964
rect 71593 1955 71651 1961
rect 71593 1921 71605 1955
rect 71639 1952 71651 1955
rect 71682 1952 71688 1964
rect 71639 1924 71688 1952
rect 71639 1921 71651 1924
rect 71593 1915 71651 1921
rect 71682 1912 71688 1924
rect 71740 1912 71746 1964
rect 73706 1912 73712 1964
rect 73764 1912 73770 1964
rect 68554 1844 68560 1896
rect 68612 1884 68618 1896
rect 69109 1887 69167 1893
rect 69109 1884 69121 1887
rect 68612 1856 69121 1884
rect 68612 1844 68618 1856
rect 69109 1853 69121 1856
rect 69155 1853 69167 1887
rect 69109 1847 69167 1853
rect 71314 1844 71320 1896
rect 71372 1884 71378 1896
rect 71869 1887 71927 1893
rect 71869 1884 71881 1887
rect 71372 1856 71881 1884
rect 71372 1844 71378 1856
rect 71869 1853 71881 1856
rect 71915 1853 71927 1887
rect 71869 1847 71927 1853
rect 70946 1816 70952 1828
rect 66732 1788 70952 1816
rect 64012 1776 64018 1788
rect 70946 1776 70952 1788
rect 71004 1776 71010 1828
rect 63862 1748 63868 1760
rect 47780 1720 63868 1748
rect 63862 1708 63868 1720
rect 63920 1708 63926 1760
rect 67450 1708 67456 1760
rect 67508 1708 67514 1760
rect 1012 1658 74980 1680
rect 1012 1606 1858 1658
rect 1910 1606 1922 1658
rect 1974 1606 1986 1658
rect 2038 1606 2050 1658
rect 2102 1606 2114 1658
rect 2166 1606 11858 1658
rect 11910 1606 11922 1658
rect 11974 1606 11986 1658
rect 12038 1606 12050 1658
rect 12102 1606 12114 1658
rect 12166 1606 21858 1658
rect 21910 1606 21922 1658
rect 21974 1606 21986 1658
rect 22038 1606 22050 1658
rect 22102 1606 22114 1658
rect 22166 1606 31858 1658
rect 31910 1606 31922 1658
rect 31974 1606 31986 1658
rect 32038 1606 32050 1658
rect 32102 1606 32114 1658
rect 32166 1606 41858 1658
rect 41910 1606 41922 1658
rect 41974 1606 41986 1658
rect 42038 1606 42050 1658
rect 42102 1606 42114 1658
rect 42166 1606 51858 1658
rect 51910 1606 51922 1658
rect 51974 1606 51986 1658
rect 52038 1606 52050 1658
rect 52102 1606 52114 1658
rect 52166 1606 61858 1658
rect 61910 1606 61922 1658
rect 61974 1606 61986 1658
rect 62038 1606 62050 1658
rect 62102 1606 62114 1658
rect 62166 1606 71858 1658
rect 71910 1606 71922 1658
rect 71974 1606 71986 1658
rect 72038 1606 72050 1658
rect 72102 1606 72114 1658
rect 72166 1606 74980 1658
rect 1012 1584 74980 1606
rect 23477 1547 23535 1553
rect 23477 1513 23489 1547
rect 23523 1544 23535 1547
rect 23566 1544 23572 1556
rect 23523 1516 23572 1544
rect 23523 1513 23535 1516
rect 23477 1507 23535 1513
rect 23566 1504 23572 1516
rect 23624 1504 23630 1556
rect 32677 1547 32735 1553
rect 32677 1513 32689 1547
rect 32723 1544 32735 1547
rect 33042 1544 33048 1556
rect 32723 1516 33048 1544
rect 32723 1513 32735 1516
rect 32677 1507 32735 1513
rect 33042 1504 33048 1516
rect 33100 1504 33106 1556
rect 35437 1547 35495 1553
rect 35437 1513 35449 1547
rect 35483 1544 35495 1547
rect 35526 1544 35532 1556
rect 35483 1516 35532 1544
rect 35483 1513 35495 1516
rect 35437 1507 35495 1513
rect 35526 1504 35532 1516
rect 35584 1504 35590 1556
rect 41322 1504 41328 1556
rect 41380 1544 41386 1556
rect 43809 1547 43867 1553
rect 43809 1544 43821 1547
rect 41380 1516 43821 1544
rect 41380 1504 41386 1516
rect 43809 1513 43821 1516
rect 43855 1513 43867 1547
rect 43809 1507 43867 1513
rect 45554 1504 45560 1556
rect 45612 1544 45618 1556
rect 46661 1547 46719 1553
rect 46661 1544 46673 1547
rect 45612 1516 46673 1544
rect 45612 1504 45618 1516
rect 46661 1513 46673 1516
rect 46707 1513 46719 1547
rect 46661 1507 46719 1513
rect 46934 1504 46940 1556
rect 46992 1544 46998 1556
rect 59722 1544 59728 1556
rect 46992 1516 59728 1544
rect 46992 1504 46998 1516
rect 59722 1504 59728 1516
rect 59780 1504 59786 1556
rect 65058 1544 65064 1556
rect 60016 1516 65064 1544
rect 21913 1479 21971 1485
rect 21913 1445 21925 1479
rect 21959 1476 21971 1479
rect 21959 1448 22692 1476
rect 21959 1445 21971 1448
rect 21913 1439 21971 1445
rect 22370 1408 22376 1420
rect 22204 1380 22376 1408
rect 20257 1343 20315 1349
rect 20257 1309 20269 1343
rect 20303 1309 20315 1343
rect 20257 1303 20315 1309
rect 20272 1272 20300 1303
rect 20990 1300 20996 1352
rect 21048 1300 21054 1352
rect 21726 1300 21732 1352
rect 21784 1300 21790 1352
rect 22005 1343 22063 1349
rect 22005 1309 22017 1343
rect 22051 1340 22063 1343
rect 22204 1340 22232 1380
rect 22370 1368 22376 1380
rect 22428 1368 22434 1420
rect 22051 1312 22232 1340
rect 22051 1309 22063 1312
rect 22005 1303 22063 1309
rect 22664 1272 22692 1448
rect 26142 1436 26148 1488
rect 26200 1476 26206 1488
rect 30834 1476 30840 1488
rect 26200 1448 30840 1476
rect 26200 1436 26206 1448
rect 30834 1436 30840 1448
rect 30892 1436 30898 1488
rect 35618 1436 35624 1488
rect 35676 1476 35682 1488
rect 60016 1476 60044 1516
rect 65058 1504 65064 1516
rect 65116 1504 65122 1556
rect 67729 1547 67787 1553
rect 67729 1513 67741 1547
rect 67775 1544 67787 1547
rect 68462 1544 68468 1556
rect 67775 1516 68468 1544
rect 67775 1513 67787 1516
rect 67729 1507 67787 1513
rect 68462 1504 68468 1516
rect 68520 1504 68526 1556
rect 73706 1504 73712 1556
rect 73764 1544 73770 1556
rect 73985 1547 74043 1553
rect 73985 1544 73997 1547
rect 73764 1516 73997 1544
rect 73764 1504 73770 1516
rect 73985 1513 73997 1516
rect 74031 1513 74043 1547
rect 73985 1507 74043 1513
rect 35676 1448 60044 1476
rect 35676 1436 35682 1448
rect 61654 1436 61660 1488
rect 61712 1476 61718 1488
rect 61841 1479 61899 1485
rect 61841 1476 61853 1479
rect 61712 1448 61853 1476
rect 61712 1436 61718 1448
rect 61841 1445 61853 1448
rect 61887 1445 61899 1479
rect 65150 1476 65156 1488
rect 61841 1439 61899 1445
rect 64846 1448 65156 1476
rect 22830 1368 22836 1420
rect 22888 1368 22894 1420
rect 32876 1380 33088 1408
rect 24121 1343 24179 1349
rect 24121 1309 24133 1343
rect 24167 1340 24179 1343
rect 25130 1340 25136 1352
rect 24167 1312 25136 1340
rect 24167 1309 24179 1312
rect 24121 1303 24179 1309
rect 25130 1300 25136 1312
rect 25188 1300 25194 1352
rect 25590 1300 25596 1352
rect 25648 1300 25654 1352
rect 26418 1300 26424 1352
rect 26476 1300 26482 1352
rect 26694 1300 26700 1352
rect 26752 1300 26758 1352
rect 27154 1300 27160 1352
rect 27212 1300 27218 1352
rect 27801 1343 27859 1349
rect 27801 1309 27813 1343
rect 27847 1340 27859 1343
rect 27847 1312 29224 1340
rect 27847 1309 27859 1312
rect 27801 1303 27859 1309
rect 20272 1244 21680 1272
rect 22664 1244 23888 1272
rect 20806 1164 20812 1216
rect 20864 1164 20870 1216
rect 21542 1164 21548 1216
rect 21600 1164 21606 1216
rect 21652 1204 21680 1244
rect 22278 1204 22284 1216
rect 21652 1176 22284 1204
rect 22278 1164 22284 1176
rect 22336 1164 22342 1216
rect 22646 1164 22652 1216
rect 22704 1164 22710 1216
rect 23382 1164 23388 1216
rect 23440 1164 23446 1216
rect 23860 1204 23888 1244
rect 23934 1232 23940 1284
rect 23992 1272 23998 1284
rect 24581 1275 24639 1281
rect 24581 1272 24593 1275
rect 23992 1244 24593 1272
rect 23992 1232 23998 1244
rect 24581 1241 24593 1244
rect 24627 1241 24639 1275
rect 24581 1235 24639 1241
rect 28353 1275 28411 1281
rect 28353 1241 28365 1275
rect 28399 1272 28411 1275
rect 28534 1272 28540 1284
rect 28399 1244 28540 1272
rect 28399 1241 28411 1244
rect 28353 1235 28411 1241
rect 28534 1232 28540 1244
rect 28592 1232 28598 1284
rect 29196 1272 29224 1312
rect 29270 1300 29276 1352
rect 29328 1300 29334 1352
rect 29825 1343 29883 1349
rect 29825 1309 29837 1343
rect 29871 1340 29883 1343
rect 29871 1312 30880 1340
rect 29871 1309 29883 1312
rect 29825 1303 29883 1309
rect 30742 1272 30748 1284
rect 29196 1244 30748 1272
rect 30742 1232 30748 1244
rect 30800 1232 30806 1284
rect 26878 1204 26884 1216
rect 23860 1176 26884 1204
rect 26878 1164 26884 1176
rect 26936 1164 26942 1216
rect 30377 1207 30435 1213
rect 30377 1173 30389 1207
rect 30423 1204 30435 1207
rect 30466 1204 30472 1216
rect 30423 1176 30472 1204
rect 30423 1173 30435 1176
rect 30377 1167 30435 1173
rect 30466 1164 30472 1176
rect 30524 1164 30530 1216
rect 30852 1204 30880 1312
rect 31570 1300 31576 1352
rect 31628 1340 31634 1352
rect 31757 1343 31815 1349
rect 31757 1340 31769 1343
rect 31628 1312 31769 1340
rect 31628 1300 31634 1312
rect 31757 1309 31769 1312
rect 31803 1309 31815 1343
rect 31757 1303 31815 1309
rect 32125 1343 32183 1349
rect 32125 1309 32137 1343
rect 32171 1340 32183 1343
rect 32876 1340 32904 1380
rect 32171 1312 32904 1340
rect 32171 1309 32183 1312
rect 32125 1303 32183 1309
rect 32950 1300 32956 1352
rect 33008 1300 33014 1352
rect 33060 1340 33088 1380
rect 38654 1368 38660 1420
rect 38712 1408 38718 1420
rect 38712 1380 41414 1408
rect 38712 1368 38718 1380
rect 34885 1343 34943 1349
rect 33060 1312 34100 1340
rect 30929 1275 30987 1281
rect 30929 1241 30941 1275
rect 30975 1272 30987 1275
rect 30975 1244 33640 1272
rect 30975 1241 30987 1244
rect 30929 1235 30987 1241
rect 33502 1204 33508 1216
rect 30852 1176 33508 1204
rect 33502 1164 33508 1176
rect 33560 1164 33566 1216
rect 33612 1204 33640 1244
rect 33962 1232 33968 1284
rect 34020 1232 34026 1284
rect 34072 1272 34100 1312
rect 34885 1309 34897 1343
rect 34931 1340 34943 1343
rect 34931 1312 36676 1340
rect 34931 1309 34943 1312
rect 34885 1303 34943 1309
rect 35066 1272 35072 1284
rect 34072 1244 35072 1272
rect 35066 1232 35072 1244
rect 35124 1232 35130 1284
rect 35434 1232 35440 1284
rect 35492 1272 35498 1284
rect 35713 1275 35771 1281
rect 35713 1272 35725 1275
rect 35492 1244 35725 1272
rect 35492 1232 35498 1244
rect 35713 1241 35725 1244
rect 35759 1241 35771 1275
rect 36538 1272 36544 1284
rect 35713 1235 35771 1241
rect 35866 1244 36544 1272
rect 35866 1204 35894 1244
rect 36538 1232 36544 1244
rect 36596 1232 36602 1284
rect 36648 1272 36676 1312
rect 36906 1300 36912 1352
rect 36964 1300 36970 1352
rect 37553 1343 37611 1349
rect 37553 1309 37565 1343
rect 37599 1340 37611 1343
rect 37599 1312 38976 1340
rect 37599 1309 37611 1312
rect 37553 1303 37611 1309
rect 37274 1272 37280 1284
rect 36648 1244 37280 1272
rect 37274 1232 37280 1244
rect 37332 1232 37338 1284
rect 38194 1232 38200 1284
rect 38252 1272 38258 1284
rect 38381 1275 38439 1281
rect 38381 1272 38393 1275
rect 38252 1244 38393 1272
rect 38252 1232 38258 1244
rect 38381 1241 38393 1244
rect 38427 1241 38439 1275
rect 38948 1272 38976 1312
rect 39390 1300 39396 1352
rect 39448 1300 39454 1352
rect 40494 1340 40500 1352
rect 39500 1312 40500 1340
rect 39500 1272 39528 1312
rect 40494 1300 40500 1312
rect 40552 1300 40558 1352
rect 41138 1300 41144 1352
rect 41196 1300 41202 1352
rect 41386 1340 41414 1380
rect 42794 1368 42800 1420
rect 42852 1408 42858 1420
rect 42852 1380 46520 1408
rect 42852 1368 42858 1380
rect 41785 1343 41843 1349
rect 41785 1340 41797 1343
rect 41386 1312 41797 1340
rect 41785 1309 41797 1312
rect 41831 1309 41843 1343
rect 41785 1303 41843 1309
rect 43717 1343 43775 1349
rect 43717 1309 43729 1343
rect 43763 1340 43775 1343
rect 43990 1340 43996 1352
rect 43763 1312 43996 1340
rect 43763 1309 43775 1312
rect 43717 1303 43775 1309
rect 43990 1300 43996 1312
rect 44048 1300 44054 1352
rect 44453 1343 44511 1349
rect 44453 1309 44465 1343
rect 44499 1340 44511 1343
rect 44818 1340 44824 1352
rect 44499 1312 44824 1340
rect 44499 1309 44511 1312
rect 44453 1303 44511 1309
rect 44818 1300 44824 1312
rect 44876 1300 44882 1352
rect 46382 1300 46388 1352
rect 46440 1300 46446 1352
rect 46492 1340 46520 1380
rect 48498 1368 48504 1420
rect 48556 1408 48562 1420
rect 49513 1411 49571 1417
rect 49513 1408 49525 1411
rect 48556 1380 49525 1408
rect 48556 1368 48562 1380
rect 49513 1377 49525 1380
rect 49559 1377 49571 1411
rect 49513 1371 49571 1377
rect 51368 1380 51580 1408
rect 47213 1343 47271 1349
rect 47213 1340 47225 1343
rect 46492 1312 47225 1340
rect 47213 1309 47225 1312
rect 47259 1309 47271 1343
rect 47213 1303 47271 1309
rect 48869 1343 48927 1349
rect 48869 1309 48881 1343
rect 48915 1340 48927 1343
rect 49050 1340 49056 1352
rect 48915 1312 49056 1340
rect 48915 1309 48927 1312
rect 48869 1303 48927 1309
rect 49050 1300 49056 1312
rect 49108 1300 49114 1352
rect 49326 1300 49332 1352
rect 49384 1340 49390 1352
rect 51368 1340 51396 1380
rect 49384 1312 51396 1340
rect 49384 1300 49390 1312
rect 51442 1300 51448 1352
rect 51500 1300 51506 1352
rect 51552 1349 51580 1380
rect 55858 1368 55864 1420
rect 55916 1408 55922 1420
rect 64846 1408 64874 1448
rect 65150 1436 65156 1448
rect 65208 1436 65214 1488
rect 55916 1380 64874 1408
rect 55916 1368 55922 1380
rect 64966 1368 64972 1420
rect 65024 1368 65030 1420
rect 67174 1368 67180 1420
rect 67232 1408 67238 1420
rect 68557 1411 68615 1417
rect 68557 1408 68569 1411
rect 67232 1380 68569 1408
rect 67232 1368 67238 1380
rect 68557 1377 68569 1380
rect 68603 1377 68615 1411
rect 68557 1371 68615 1377
rect 69934 1368 69940 1420
rect 69992 1408 69998 1420
rect 71133 1411 71191 1417
rect 71133 1408 71145 1411
rect 69992 1380 71145 1408
rect 69992 1368 69998 1380
rect 71133 1377 71145 1380
rect 71179 1377 71191 1411
rect 71133 1371 71191 1377
rect 74626 1368 74632 1420
rect 74684 1368 74690 1420
rect 51537 1343 51595 1349
rect 51537 1309 51549 1343
rect 51583 1309 51595 1343
rect 51537 1303 51595 1309
rect 51626 1300 51632 1352
rect 51684 1340 51690 1352
rect 52089 1343 52147 1349
rect 52089 1340 52101 1343
rect 51684 1312 52101 1340
rect 51684 1300 51690 1312
rect 52089 1309 52101 1312
rect 52135 1309 52147 1343
rect 52089 1303 52147 1309
rect 54018 1300 54024 1352
rect 54076 1300 54082 1352
rect 54665 1343 54723 1349
rect 54665 1309 54677 1343
rect 54711 1309 54723 1343
rect 54665 1303 54723 1309
rect 56505 1343 56563 1349
rect 56505 1309 56517 1343
rect 56551 1309 56563 1343
rect 56505 1303 56563 1309
rect 38948 1244 39528 1272
rect 38381 1235 38439 1241
rect 39574 1232 39580 1284
rect 39632 1272 39638 1284
rect 40037 1275 40095 1281
rect 40037 1272 40049 1275
rect 39632 1244 40049 1272
rect 39632 1232 39638 1244
rect 40037 1241 40049 1244
rect 40083 1241 40095 1275
rect 40037 1235 40095 1241
rect 40126 1232 40132 1284
rect 40184 1272 40190 1284
rect 41233 1275 41291 1281
rect 41233 1272 41245 1275
rect 40184 1244 41245 1272
rect 40184 1232 40190 1244
rect 41233 1241 41245 1244
rect 41279 1241 41291 1275
rect 41233 1235 41291 1241
rect 41322 1232 41328 1284
rect 41380 1272 41386 1284
rect 42521 1275 42579 1281
rect 42521 1272 42533 1275
rect 41380 1244 42533 1272
rect 41380 1232 41386 1244
rect 42521 1241 42533 1244
rect 42567 1241 42579 1275
rect 42521 1235 42579 1241
rect 45094 1232 45100 1284
rect 45152 1272 45158 1284
rect 45373 1275 45431 1281
rect 45373 1272 45385 1275
rect 45152 1244 45385 1272
rect 45152 1232 45158 1244
rect 45373 1241 45385 1244
rect 45419 1241 45431 1275
rect 45373 1235 45431 1241
rect 46474 1232 46480 1284
rect 46532 1272 46538 1284
rect 47673 1275 47731 1281
rect 47673 1272 47685 1275
rect 46532 1244 47685 1272
rect 46532 1232 46538 1244
rect 47673 1241 47685 1244
rect 47719 1241 47731 1275
rect 47673 1235 47731 1241
rect 48314 1232 48320 1284
rect 48372 1272 48378 1284
rect 48961 1275 49019 1281
rect 48961 1272 48973 1275
rect 48372 1244 48973 1272
rect 48372 1232 48378 1244
rect 48961 1241 48973 1244
rect 49007 1241 49019 1275
rect 48961 1235 49019 1241
rect 49234 1232 49240 1284
rect 49292 1272 49298 1284
rect 50249 1275 50307 1281
rect 50249 1272 50261 1275
rect 49292 1244 50261 1272
rect 49292 1232 49298 1244
rect 50249 1241 50261 1244
rect 50295 1241 50307 1275
rect 50249 1235 50307 1241
rect 51046 1244 51672 1272
rect 33612 1176 35894 1204
rect 38105 1207 38163 1213
rect 38105 1173 38117 1207
rect 38151 1204 38163 1207
rect 41046 1204 41052 1216
rect 38151 1176 41052 1204
rect 38151 1173 38163 1176
rect 38105 1167 38163 1173
rect 41046 1164 41052 1176
rect 41104 1164 41110 1216
rect 50154 1164 50160 1216
rect 50212 1204 50218 1216
rect 51046 1204 51074 1244
rect 50212 1176 51074 1204
rect 51644 1204 51672 1244
rect 52362 1232 52368 1284
rect 52420 1272 52426 1284
rect 52825 1275 52883 1281
rect 52825 1272 52837 1275
rect 52420 1244 52837 1272
rect 52420 1232 52426 1244
rect 52825 1241 52837 1244
rect 52871 1241 52883 1275
rect 54680 1272 54708 1303
rect 52825 1235 52883 1241
rect 52932 1244 54708 1272
rect 52932 1204 52960 1244
rect 54754 1232 54760 1284
rect 54812 1272 54818 1284
rect 55401 1275 55459 1281
rect 55401 1272 55413 1275
rect 54812 1244 55413 1272
rect 54812 1232 54818 1244
rect 55401 1241 55413 1244
rect 55447 1241 55459 1275
rect 55401 1235 55459 1241
rect 51644 1176 52960 1204
rect 50212 1164 50218 1176
rect 53926 1164 53932 1216
rect 53984 1204 53990 1216
rect 54113 1207 54171 1213
rect 54113 1204 54125 1207
rect 53984 1176 54125 1204
rect 53984 1164 53990 1176
rect 54113 1173 54125 1176
rect 54159 1173 54171 1207
rect 56520 1204 56548 1303
rect 56686 1300 56692 1352
rect 56744 1300 56750 1352
rect 57238 1300 57244 1352
rect 57296 1300 57302 1352
rect 59078 1300 59084 1352
rect 59136 1300 59142 1352
rect 59262 1300 59268 1352
rect 59320 1300 59326 1352
rect 59446 1300 59452 1352
rect 59504 1340 59510 1352
rect 59817 1343 59875 1349
rect 59817 1340 59829 1343
rect 59504 1312 59829 1340
rect 59504 1300 59510 1312
rect 59817 1309 59829 1312
rect 59863 1309 59875 1343
rect 59817 1303 59875 1309
rect 61749 1343 61807 1349
rect 61749 1309 61761 1343
rect 61795 1340 61807 1343
rect 62298 1340 62304 1352
rect 61795 1312 62304 1340
rect 61795 1309 61807 1312
rect 61749 1303 61807 1309
rect 62298 1300 62304 1312
rect 62356 1300 62362 1352
rect 62390 1300 62396 1352
rect 62448 1300 62454 1352
rect 63126 1300 63132 1352
rect 63184 1300 63190 1352
rect 63402 1300 63408 1352
rect 63460 1340 63466 1352
rect 64417 1343 64475 1349
rect 64417 1340 64429 1343
rect 63460 1312 64429 1340
rect 63460 1300 63466 1312
rect 64417 1309 64429 1312
rect 64463 1309 64475 1343
rect 64417 1303 64475 1309
rect 65886 1300 65892 1352
rect 65944 1300 65950 1352
rect 67450 1300 67456 1352
rect 67508 1300 67514 1352
rect 68186 1300 68192 1352
rect 68244 1300 68250 1352
rect 69382 1300 69388 1352
rect 69440 1340 69446 1352
rect 69569 1343 69627 1349
rect 69569 1340 69581 1343
rect 69440 1312 69581 1340
rect 69440 1300 69446 1312
rect 69569 1309 69581 1312
rect 69615 1309 69627 1343
rect 69569 1303 69627 1309
rect 69750 1300 69756 1352
rect 69808 1340 69814 1352
rect 70121 1343 70179 1349
rect 70121 1340 70133 1343
rect 69808 1312 70133 1340
rect 69808 1300 69814 1312
rect 70121 1309 70133 1312
rect 70167 1309 70179 1343
rect 70121 1303 70179 1309
rect 70762 1300 70768 1352
rect 70820 1300 70826 1352
rect 72145 1343 72203 1349
rect 72145 1309 72157 1343
rect 72191 1340 72203 1343
rect 72234 1340 72240 1352
rect 72191 1312 72240 1340
rect 72191 1309 72203 1312
rect 72145 1303 72203 1309
rect 72234 1300 72240 1312
rect 72292 1300 72298 1352
rect 72694 1300 72700 1352
rect 72752 1300 72758 1352
rect 73246 1300 73252 1352
rect 73304 1300 73310 1352
rect 73801 1343 73859 1349
rect 73801 1309 73813 1343
rect 73847 1309 73859 1343
rect 73801 1303 73859 1309
rect 57514 1232 57520 1284
rect 57572 1272 57578 1284
rect 57977 1275 58035 1281
rect 57977 1272 57989 1275
rect 57572 1244 57989 1272
rect 57572 1232 57578 1244
rect 57977 1241 57989 1244
rect 58023 1241 58035 1275
rect 57977 1235 58035 1241
rect 60274 1232 60280 1284
rect 60332 1272 60338 1284
rect 60553 1275 60611 1281
rect 60553 1272 60565 1275
rect 60332 1244 60565 1272
rect 60332 1232 60338 1244
rect 60553 1241 60565 1244
rect 60599 1241 60611 1275
rect 60553 1235 60611 1241
rect 61654 1232 61660 1284
rect 61712 1272 61718 1284
rect 63865 1275 63923 1281
rect 63865 1272 63877 1275
rect 61712 1244 63877 1272
rect 61712 1232 61718 1244
rect 63865 1241 63877 1244
rect 63911 1241 63923 1275
rect 63865 1235 63923 1241
rect 65794 1232 65800 1284
rect 65852 1272 65858 1284
rect 66809 1275 66867 1281
rect 66809 1272 66821 1275
rect 65852 1244 66821 1272
rect 65852 1232 65858 1244
rect 66809 1241 66821 1244
rect 66855 1241 66867 1275
rect 66809 1235 66867 1241
rect 70854 1232 70860 1284
rect 70912 1272 70918 1284
rect 73816 1272 73844 1303
rect 70912 1244 73844 1272
rect 70912 1232 70918 1244
rect 63678 1204 63684 1216
rect 56520 1176 63684 1204
rect 54113 1167 54171 1173
rect 63678 1164 63684 1176
rect 63736 1164 63742 1216
rect 1012 1114 74980 1136
rect 1012 1062 4210 1114
rect 4262 1062 4274 1114
rect 4326 1062 4338 1114
rect 4390 1062 4402 1114
rect 4454 1062 4466 1114
rect 4518 1062 14210 1114
rect 14262 1062 14274 1114
rect 14326 1062 14338 1114
rect 14390 1062 14402 1114
rect 14454 1062 14466 1114
rect 14518 1062 24210 1114
rect 24262 1062 24274 1114
rect 24326 1062 24338 1114
rect 24390 1062 24402 1114
rect 24454 1062 24466 1114
rect 24518 1062 34210 1114
rect 34262 1062 34274 1114
rect 34326 1062 34338 1114
rect 34390 1062 34402 1114
rect 34454 1062 34466 1114
rect 34518 1062 44210 1114
rect 44262 1062 44274 1114
rect 44326 1062 44338 1114
rect 44390 1062 44402 1114
rect 44454 1062 44466 1114
rect 44518 1062 54210 1114
rect 54262 1062 54274 1114
rect 54326 1062 54338 1114
rect 54390 1062 54402 1114
rect 54454 1062 54466 1114
rect 54518 1062 64210 1114
rect 64262 1062 64274 1114
rect 64326 1062 64338 1114
rect 64390 1062 64402 1114
rect 64454 1062 64466 1114
rect 64518 1062 74210 1114
rect 74262 1062 74274 1114
rect 74326 1062 74338 1114
rect 74390 1062 74402 1114
rect 74454 1062 74466 1114
rect 74518 1062 74980 1114
rect 1012 1040 74980 1062
rect 21726 960 21732 1012
rect 21784 1000 21790 1012
rect 23290 1000 23296 1012
rect 21784 972 23296 1000
rect 21784 960 21790 972
rect 23290 960 23296 972
rect 23348 960 23354 1012
rect 23382 960 23388 1012
rect 23440 1000 23446 1012
rect 26510 1000 26516 1012
rect 23440 972 26516 1000
rect 23440 960 23446 972
rect 26510 960 26516 972
rect 26568 960 26574 1012
rect 30466 960 30472 1012
rect 30524 1000 30530 1012
rect 33870 1000 33876 1012
rect 30524 972 33876 1000
rect 30524 960 30530 972
rect 33870 960 33876 972
rect 33928 960 33934 1012
rect 36538 960 36544 1012
rect 36596 1000 36602 1012
rect 39758 1000 39764 1012
rect 36596 972 39764 1000
rect 36596 960 36602 972
rect 39758 960 39764 972
rect 39816 960 39822 1012
rect 41138 960 41144 1012
rect 41196 1000 41202 1012
rect 65978 1000 65984 1012
rect 41196 972 65984 1000
rect 41196 960 41202 972
rect 65978 960 65984 972
rect 66036 960 66042 1012
rect 20806 892 20812 944
rect 20864 932 20870 944
rect 23658 932 23664 944
rect 20864 904 23664 932
rect 20864 892 20870 904
rect 23658 892 23664 904
rect 23716 892 23722 944
rect 28994 892 29000 944
rect 29052 892 29058 944
rect 33962 892 33968 944
rect 34020 932 34026 944
rect 40402 932 40408 944
rect 34020 904 40408 932
rect 34020 892 34026 904
rect 40402 892 40408 904
rect 40460 892 40466 944
rect 49050 892 49056 944
rect 49108 932 49114 944
rect 72602 932 72608 944
rect 49108 904 72608 932
rect 49108 892 49114 904
rect 72602 892 72608 904
rect 72660 892 72666 944
rect 22370 824 22376 876
rect 22428 864 22434 876
rect 26050 864 26056 876
rect 22428 836 26056 864
rect 22428 824 22434 836
rect 26050 824 26056 836
rect 26108 824 26114 876
rect 21542 756 21548 808
rect 21600 796 21606 808
rect 25038 796 25044 808
rect 21600 768 25044 796
rect 21600 756 21606 768
rect 25038 756 25044 768
rect 25096 756 25102 808
rect 25130 756 25136 808
rect 25188 796 25194 808
rect 29012 796 29040 892
rect 43990 824 43996 876
rect 44048 864 44054 876
rect 65426 864 65432 876
rect 44048 836 65432 864
rect 44048 824 44054 836
rect 65426 824 65432 836
rect 65484 824 65490 876
rect 25188 768 29040 796
rect 25188 756 25194 768
rect 29270 756 29276 808
rect 29328 796 29334 808
rect 64046 796 64052 808
rect 29328 768 64052 796
rect 29328 756 29334 768
rect 64046 756 64052 768
rect 64104 756 64110 808
rect 22646 688 22652 740
rect 22704 728 22710 740
rect 28350 728 28356 740
rect 22704 700 28356 728
rect 22704 688 22710 700
rect 28350 688 28356 700
rect 28408 688 28414 740
rect 46382 688 46388 740
rect 46440 728 46446 740
rect 70486 728 70492 740
rect 46440 700 70492 728
rect 46440 688 46446 700
rect 70486 688 70492 700
rect 70544 688 70550 740
rect 36906 620 36912 672
rect 36964 660 36970 672
rect 65242 660 65248 672
rect 36964 632 65248 660
rect 36964 620 36970 632
rect 65242 620 65248 632
rect 65300 620 65306 672
rect 39390 552 39396 604
rect 39448 592 39454 604
rect 64966 592 64972 604
rect 39448 564 64972 592
rect 39448 552 39454 564
rect 64966 552 64972 564
rect 65024 552 65030 604
rect 54018 484 54024 536
rect 54076 524 54082 536
rect 63770 524 63776 536
rect 54076 496 63776 524
rect 54076 484 54082 496
rect 63770 484 63776 496
rect 63828 484 63834 536
rect 63126 348 63132 400
rect 63184 388 63190 400
rect 72786 388 72792 400
rect 63184 360 72792 388
rect 63184 348 63190 360
rect 72786 348 72792 360
rect 72844 348 72850 400
rect 51442 280 51448 332
rect 51500 320 51506 332
rect 65610 320 65616 332
rect 51500 292 65616 320
rect 51500 280 51506 292
rect 65610 280 65616 292
rect 65668 280 65674 332
<< via1 >>
rect 74210 85926 74262 85978
rect 74274 85926 74326 85978
rect 74338 85926 74390 85978
rect 74402 85926 74454 85978
rect 74466 85926 74518 85978
rect 71858 85382 71910 85434
rect 71922 85382 71974 85434
rect 71986 85382 72038 85434
rect 72050 85382 72102 85434
rect 72114 85382 72166 85434
rect 74210 84838 74262 84890
rect 74274 84838 74326 84890
rect 74338 84838 74390 84890
rect 74402 84838 74454 84890
rect 74466 84838 74518 84890
rect 71858 84294 71910 84346
rect 71922 84294 71974 84346
rect 71986 84294 72038 84346
rect 72050 84294 72102 84346
rect 72114 84294 72166 84346
rect 64880 84192 64932 84244
rect 74210 83750 74262 83802
rect 74274 83750 74326 83802
rect 74338 83750 74390 83802
rect 74402 83750 74454 83802
rect 74466 83750 74518 83802
rect 71858 83206 71910 83258
rect 71922 83206 71974 83258
rect 71986 83206 72038 83258
rect 72050 83206 72102 83258
rect 72114 83206 72166 83258
rect 65708 83104 65760 83156
rect 71688 82968 71740 83020
rect 74210 82662 74262 82714
rect 74274 82662 74326 82714
rect 74338 82662 74390 82714
rect 74402 82662 74454 82714
rect 74466 82662 74518 82714
rect 71858 82118 71910 82170
rect 71922 82118 71974 82170
rect 71986 82118 72038 82170
rect 72050 82118 72102 82170
rect 72114 82118 72166 82170
rect 64880 81744 64932 81796
rect 74210 81574 74262 81626
rect 74274 81574 74326 81626
rect 74338 81574 74390 81626
rect 74402 81574 74454 81626
rect 74466 81574 74518 81626
rect 71858 81030 71910 81082
rect 71922 81030 71974 81082
rect 71986 81030 72038 81082
rect 72050 81030 72102 81082
rect 72114 81030 72166 81082
rect 65524 80928 65576 80980
rect 70676 80792 70728 80844
rect 74210 80486 74262 80538
rect 74274 80486 74326 80538
rect 74338 80486 74390 80538
rect 74402 80486 74454 80538
rect 74466 80486 74518 80538
rect 71858 79942 71910 79994
rect 71922 79942 71974 79994
rect 71986 79942 72038 79994
rect 72050 79942 72102 79994
rect 72114 79942 72166 79994
rect 64880 79840 64932 79892
rect 74210 79398 74262 79450
rect 74274 79398 74326 79450
rect 74338 79398 74390 79450
rect 74402 79398 74454 79450
rect 74466 79398 74518 79450
rect 71858 78854 71910 78906
rect 71922 78854 71974 78906
rect 71986 78854 72038 78906
rect 72050 78854 72102 78906
rect 72114 78854 72166 78906
rect 65616 78684 65668 78736
rect 68652 78616 68704 78668
rect 74210 78310 74262 78362
rect 74274 78310 74326 78362
rect 74338 78310 74390 78362
rect 74402 78310 74454 78362
rect 74466 78310 74518 78362
rect 71858 77766 71910 77818
rect 71922 77766 71974 77818
rect 71986 77766 72038 77818
rect 72050 77766 72102 77818
rect 72114 77766 72166 77818
rect 64880 77664 64932 77716
rect 74210 77222 74262 77274
rect 74274 77222 74326 77274
rect 74338 77222 74390 77274
rect 74402 77222 74454 77274
rect 74466 77222 74518 77274
rect 71858 76678 71910 76730
rect 71922 76678 71974 76730
rect 71986 76678 72038 76730
rect 72050 76678 72102 76730
rect 72114 76678 72166 76730
rect 65340 76508 65392 76560
rect 68100 76440 68152 76492
rect 74210 76134 74262 76186
rect 74274 76134 74326 76186
rect 74338 76134 74390 76186
rect 74402 76134 74454 76186
rect 74466 76134 74518 76186
rect 71858 75590 71910 75642
rect 71922 75590 71974 75642
rect 71986 75590 72038 75642
rect 72050 75590 72102 75642
rect 72114 75590 72166 75642
rect 64880 75148 64932 75200
rect 74210 75046 74262 75098
rect 74274 75046 74326 75098
rect 74338 75046 74390 75098
rect 74402 75046 74454 75098
rect 74466 75046 74518 75098
rect 65432 74604 65484 74656
rect 71858 74502 71910 74554
rect 71922 74502 71974 74554
rect 71986 74502 72038 74554
rect 72050 74502 72102 74554
rect 72114 74502 72166 74554
rect 65892 74060 65944 74112
rect 74210 73958 74262 74010
rect 74274 73958 74326 74010
rect 74338 73958 74390 74010
rect 74402 73958 74454 74010
rect 74466 73958 74518 74010
rect 71858 73414 71910 73466
rect 71922 73414 71974 73466
rect 71986 73414 72038 73466
rect 72050 73414 72102 73466
rect 72114 73414 72166 73466
rect 64880 73176 64932 73228
rect 74210 72870 74262 72922
rect 74274 72870 74326 72922
rect 74338 72870 74390 72922
rect 74402 72870 74454 72922
rect 74466 72870 74518 72922
rect 71858 72326 71910 72378
rect 71922 72326 71974 72378
rect 71986 72326 72038 72378
rect 72050 72326 72102 72378
rect 72114 72326 72166 72378
rect 65156 72156 65208 72208
rect 64604 71748 64656 71800
rect 74210 71782 74262 71834
rect 74274 71782 74326 71834
rect 74338 71782 74390 71834
rect 74402 71782 74454 71834
rect 74466 71782 74518 71834
rect 71858 71238 71910 71290
rect 71922 71238 71974 71290
rect 71986 71238 72038 71290
rect 72050 71238 72102 71290
rect 72114 71238 72166 71290
rect 64880 71068 64932 71120
rect 74210 70694 74262 70746
rect 74274 70694 74326 70746
rect 74338 70694 74390 70746
rect 74402 70694 74454 70746
rect 74466 70694 74518 70746
rect 71858 70150 71910 70202
rect 71922 70150 71974 70202
rect 71986 70150 72038 70202
rect 72050 70150 72102 70202
rect 72114 70150 72166 70202
rect 65248 69980 65300 70032
rect 71136 69912 71188 69964
rect 74210 69606 74262 69658
rect 74274 69606 74326 69658
rect 74338 69606 74390 69658
rect 74402 69606 74454 69658
rect 74466 69606 74518 69658
rect 71858 69062 71910 69114
rect 71922 69062 71974 69114
rect 71986 69062 72038 69114
rect 72050 69062 72102 69114
rect 72114 69062 72166 69114
rect 64880 68892 64932 68944
rect 65800 68892 65852 68944
rect 74210 68518 74262 68570
rect 74274 68518 74326 68570
rect 74338 68518 74390 68570
rect 74402 68518 74454 68570
rect 74466 68518 74518 68570
rect 71858 67974 71910 68026
rect 71922 67974 71974 68026
rect 71986 67974 72038 68026
rect 72050 67974 72102 68026
rect 72114 67974 72166 68026
rect 65064 67804 65116 67856
rect 72792 67736 72844 67788
rect 74210 67430 74262 67482
rect 74274 67430 74326 67482
rect 74338 67430 74390 67482
rect 74402 67430 74454 67482
rect 74466 67430 74518 67482
rect 71858 66886 71910 66938
rect 71922 66886 71974 66938
rect 71986 66886 72038 66938
rect 72050 66886 72102 66938
rect 72114 66886 72166 66938
rect 64880 66444 64932 66496
rect 74210 66342 74262 66394
rect 74274 66342 74326 66394
rect 74338 66342 74390 66394
rect 74402 66342 74454 66394
rect 74466 66342 74518 66394
rect 71858 65798 71910 65850
rect 71922 65798 71974 65850
rect 71986 65798 72038 65850
rect 72050 65798 72102 65850
rect 72114 65798 72166 65850
rect 65984 65628 66036 65680
rect 66076 65356 66128 65408
rect 74210 65254 74262 65306
rect 74274 65254 74326 65306
rect 74338 65254 74390 65306
rect 74402 65254 74454 65306
rect 74466 65254 74518 65306
rect 71858 64710 71910 64762
rect 71922 64710 71974 64762
rect 71986 64710 72038 64762
rect 72050 64710 72102 64762
rect 72114 64710 72166 64762
rect 64880 64268 64932 64320
rect 74210 64166 74262 64218
rect 74274 64166 74326 64218
rect 74338 64166 74390 64218
rect 74402 64166 74454 64218
rect 74466 64166 74518 64218
rect 71858 63622 71910 63674
rect 71922 63622 71974 63674
rect 71986 63622 72038 63674
rect 72050 63622 72102 63674
rect 72114 63622 72166 63674
rect 64972 63520 65024 63572
rect 65708 63495 65760 63504
rect 65708 63461 65717 63495
rect 65717 63461 65751 63495
rect 65751 63461 65760 63495
rect 65708 63452 65760 63461
rect 68008 63316 68060 63368
rect 63592 63044 63644 63096
rect 74210 63078 74262 63130
rect 74274 63078 74326 63130
rect 74338 63078 74390 63130
rect 74402 63078 74454 63130
rect 74466 63078 74518 63130
rect 71858 62534 71910 62586
rect 71922 62534 71974 62586
rect 71986 62534 72038 62586
rect 72050 62534 72102 62586
rect 72114 62534 72166 62586
rect 64880 62092 64932 62144
rect 74210 61990 74262 62042
rect 74274 61990 74326 62042
rect 74338 61990 74390 62042
rect 74402 61990 74454 62042
rect 74466 61990 74518 62042
rect 65524 61888 65576 61940
rect 66536 61684 66588 61736
rect 71858 61446 71910 61498
rect 71922 61446 71974 61498
rect 71986 61446 72038 61498
rect 72050 61446 72102 61498
rect 72114 61446 72166 61498
rect 66168 61276 66220 61328
rect 63500 61178 63552 61230
rect 74210 60902 74262 60954
rect 74274 60902 74326 60954
rect 74338 60902 74390 60954
rect 74402 60902 74454 60954
rect 74466 60902 74518 60954
rect 71858 60358 71910 60410
rect 71922 60358 71974 60410
rect 71986 60358 72038 60410
rect 72050 60358 72102 60410
rect 72114 60358 72166 60410
rect 65616 60299 65668 60308
rect 65616 60265 65625 60299
rect 65625 60265 65659 60299
rect 65659 60265 65668 60299
rect 65616 60256 65668 60265
rect 64880 60188 64932 60240
rect 67088 60052 67140 60104
rect 74210 59814 74262 59866
rect 74274 59814 74326 59866
rect 74338 59814 74390 59866
rect 74402 59814 74454 59866
rect 74466 59814 74518 59866
rect 71858 59270 71910 59322
rect 71922 59270 71974 59322
rect 71986 59270 72038 59322
rect 72050 59270 72102 59322
rect 72114 59270 72166 59322
rect 65708 59100 65760 59152
rect 71320 59032 71372 59084
rect 74210 58726 74262 58778
rect 74274 58726 74326 58778
rect 74338 58726 74390 58778
rect 74402 58726 74454 58778
rect 74466 58726 74518 58778
rect 65340 58624 65392 58676
rect 66260 58463 66312 58472
rect 66260 58429 66269 58463
rect 66269 58429 66303 58463
rect 66303 58429 66312 58463
rect 66260 58420 66312 58429
rect 71858 58182 71910 58234
rect 71922 58182 71974 58234
rect 71986 58182 72038 58234
rect 72050 58182 72102 58234
rect 72114 58182 72166 58234
rect 64880 58012 64932 58064
rect 74210 57638 74262 57690
rect 74274 57638 74326 57690
rect 74338 57638 74390 57690
rect 74402 57638 74454 57690
rect 74466 57638 74518 57690
rect 71858 57094 71910 57146
rect 71922 57094 71974 57146
rect 71986 57094 72038 57146
rect 72050 57094 72102 57146
rect 72114 57094 72166 57146
rect 65432 56992 65484 57044
rect 65524 56924 65576 56976
rect 69296 56788 69348 56840
rect 63684 56584 63736 56636
rect 74210 56550 74262 56602
rect 74274 56550 74326 56602
rect 74338 56550 74390 56602
rect 74402 56550 74454 56602
rect 74466 56550 74518 56602
rect 71858 56006 71910 56058
rect 71922 56006 71974 56058
rect 71986 56006 72038 56058
rect 72050 56006 72102 56058
rect 72114 56006 72166 56058
rect 64880 55564 64932 55616
rect 74210 55462 74262 55514
rect 74274 55462 74326 55514
rect 74338 55462 74390 55514
rect 74402 55462 74454 55514
rect 74466 55462 74518 55514
rect 65156 55360 65208 55412
rect 69112 55224 69164 55276
rect 71858 54918 71910 54970
rect 71922 54918 71974 54970
rect 71986 54918 72038 54970
rect 72050 54918 72102 54970
rect 72114 54918 72166 54970
rect 65340 54748 65392 54800
rect 71228 54612 71280 54664
rect 74210 54374 74262 54426
rect 74274 54374 74326 54426
rect 74338 54374 74390 54426
rect 74402 54374 74454 54426
rect 74466 54374 74518 54426
rect 71858 53830 71910 53882
rect 71922 53830 71974 53882
rect 71986 53830 72038 53882
rect 72050 53830 72102 53882
rect 72114 53830 72166 53882
rect 65800 53635 65852 53644
rect 65800 53601 65809 53635
rect 65809 53601 65843 53635
rect 65843 53601 65852 53635
rect 65800 53592 65852 53601
rect 64880 53524 64932 53576
rect 69388 53524 69440 53576
rect 69020 53388 69072 53440
rect 74210 53286 74262 53338
rect 74274 53286 74326 53338
rect 74338 53286 74390 53338
rect 74402 53286 74454 53338
rect 74466 53286 74518 53338
rect 65248 53184 65300 53236
rect 66352 52980 66404 53032
rect 71858 52742 71910 52794
rect 71922 52742 71974 52794
rect 71986 52742 72038 52794
rect 72050 52742 72102 52794
rect 72114 52742 72166 52794
rect 65432 52572 65484 52624
rect 63776 52436 63828 52488
rect 65616 52479 65668 52488
rect 65616 52445 65625 52479
rect 65625 52445 65659 52479
rect 65659 52445 65668 52479
rect 65616 52436 65668 52445
rect 74210 52198 74262 52250
rect 74274 52198 74326 52250
rect 74338 52198 74390 52250
rect 74402 52198 74454 52250
rect 74466 52198 74518 52250
rect 65616 52096 65668 52148
rect 65064 51960 65116 52012
rect 67548 51892 67600 51944
rect 71858 51654 71910 51706
rect 71922 51654 71974 51706
rect 71986 51654 72038 51706
rect 72050 51654 72102 51706
rect 72114 51654 72166 51706
rect 64880 51484 64932 51536
rect 65800 51484 65852 51536
rect 74210 51110 74262 51162
rect 74274 51110 74326 51162
rect 74338 51110 74390 51162
rect 74402 51110 74454 51162
rect 74466 51110 74518 51162
rect 71858 50566 71910 50618
rect 71922 50566 71974 50618
rect 71986 50566 72038 50618
rect 72050 50566 72102 50618
rect 72114 50566 72166 50618
rect 65984 50464 66036 50516
rect 65156 50396 65208 50448
rect 67640 50328 67692 50380
rect 63868 50260 63920 50312
rect 74210 50022 74262 50074
rect 74274 50022 74326 50074
rect 74338 50022 74390 50074
rect 74402 50022 74454 50074
rect 74466 50022 74518 50074
rect 71858 49478 71910 49530
rect 71922 49478 71974 49530
rect 71986 49478 72038 49530
rect 72050 49478 72102 49530
rect 72114 49478 72166 49530
rect 63408 49172 63460 49224
rect 74210 48934 74262 48986
rect 74274 48934 74326 48986
rect 74338 48934 74390 48986
rect 74402 48934 74454 48986
rect 74466 48934 74518 48986
rect 64972 48832 65024 48884
rect 69756 48764 69808 48816
rect 63408 48689 63460 48741
rect 69572 48628 69624 48680
rect 71858 48390 71910 48442
rect 71922 48390 71974 48442
rect 71986 48390 72038 48442
rect 72050 48390 72102 48442
rect 72114 48390 72166 48442
rect 69204 48084 69256 48136
rect 74210 47846 74262 47898
rect 74274 47846 74326 47898
rect 74338 47846 74390 47898
rect 74402 47846 74454 47898
rect 74466 47846 74518 47898
rect 64972 47676 65024 47728
rect 64880 47336 64932 47388
rect 63408 47273 63460 47325
rect 71858 47302 71910 47354
rect 71922 47302 71974 47354
rect 71986 47302 72038 47354
rect 72050 47302 72102 47354
rect 72114 47302 72166 47354
rect 66168 47200 66220 47252
rect 70768 47064 70820 47116
rect 69664 46996 69716 47048
rect 66628 46971 66680 46980
rect 66628 46937 66637 46971
rect 66637 46937 66671 46971
rect 66671 46937 66680 46971
rect 66628 46928 66680 46937
rect 74210 46758 74262 46810
rect 74274 46758 74326 46810
rect 74338 46758 74390 46810
rect 74402 46758 74454 46810
rect 74466 46758 74518 46810
rect 71858 46214 71910 46266
rect 71922 46214 71974 46266
rect 71986 46214 72038 46266
rect 72050 46214 72102 46266
rect 72114 46214 72166 46266
rect 65064 45908 65116 45960
rect 74210 45670 74262 45722
rect 74274 45670 74326 45722
rect 74338 45670 74390 45722
rect 74402 45670 74454 45722
rect 74466 45670 74518 45722
rect 66996 45568 67048 45620
rect 65616 45543 65668 45552
rect 65616 45509 65625 45543
rect 65625 45509 65659 45543
rect 65659 45509 65668 45543
rect 65616 45500 65668 45509
rect 67180 45364 67232 45416
rect 67272 45228 67324 45280
rect 71858 45126 71910 45178
rect 71922 45126 71974 45178
rect 71986 45126 72038 45178
rect 72050 45126 72102 45178
rect 72114 45126 72166 45178
rect 66812 44820 66864 44872
rect 64972 44684 65024 44736
rect 65616 44684 65668 44736
rect 64972 44548 65024 44600
rect 74210 44582 74262 44634
rect 74274 44582 74326 44634
rect 74338 44582 74390 44634
rect 74402 44582 74454 44634
rect 74466 44582 74518 44634
rect 65800 44140 65852 44192
rect 66628 44140 66680 44192
rect 70860 44140 70912 44192
rect 71858 44038 71910 44090
rect 71922 44038 71974 44090
rect 71986 44038 72038 44090
rect 72050 44038 72102 44090
rect 72114 44038 72166 44090
rect 65524 43936 65576 43988
rect 66444 43800 66496 43852
rect 65984 43732 66036 43784
rect 74210 43494 74262 43546
rect 74274 43494 74326 43546
rect 74338 43494 74390 43546
rect 74402 43494 74454 43546
rect 74466 43494 74518 43546
rect 63960 43120 64012 43172
rect 71858 42950 71910 43002
rect 71922 42950 71974 43002
rect 71986 42950 72038 43002
rect 72050 42950 72102 43002
rect 72114 42950 72166 43002
rect 66168 42780 66220 42832
rect 68008 42755 68060 42764
rect 68008 42721 68017 42755
rect 68017 42721 68051 42755
rect 68051 42721 68060 42755
rect 68008 42712 68060 42721
rect 70124 42644 70176 42696
rect 74210 42406 74262 42458
rect 74274 42406 74326 42458
rect 74338 42406 74390 42458
rect 74402 42406 74454 42458
rect 74466 42406 74518 42458
rect 65340 42304 65392 42356
rect 66720 42100 66772 42152
rect 65432 42032 65484 42084
rect 71858 41862 71910 41914
rect 71922 41862 71974 41914
rect 71986 41862 72038 41914
rect 72050 41862 72102 41914
rect 72114 41862 72166 41914
rect 65432 41760 65484 41812
rect 66536 41760 66588 41812
rect 65156 41692 65208 41744
rect 68560 41556 68612 41608
rect 74210 41318 74262 41370
rect 74274 41318 74326 41370
rect 74338 41318 74390 41370
rect 74402 41318 74454 41370
rect 74466 41318 74518 41370
rect 64052 40944 64104 40996
rect 65800 40919 65852 40928
rect 65800 40885 65809 40919
rect 65809 40885 65843 40919
rect 65843 40885 65852 40919
rect 65800 40876 65852 40885
rect 71858 40774 71910 40826
rect 71922 40774 71974 40826
rect 71986 40774 72038 40826
rect 72050 40774 72102 40826
rect 72114 40774 72166 40826
rect 67088 40715 67140 40724
rect 67088 40681 67097 40715
rect 67097 40681 67131 40715
rect 67131 40681 67140 40715
rect 67088 40672 67140 40681
rect 65340 40536 65392 40588
rect 65708 40536 65760 40588
rect 66536 40468 66588 40520
rect 68192 40468 68244 40520
rect 65708 40332 65760 40384
rect 65984 40332 66036 40384
rect 74210 40230 74262 40282
rect 74274 40230 74326 40282
rect 74338 40230 74390 40282
rect 74402 40230 74454 40282
rect 74466 40230 74518 40282
rect 65432 40128 65484 40180
rect 66628 39924 66680 39976
rect 65156 39788 65208 39840
rect 71858 39686 71910 39738
rect 71922 39686 71974 39738
rect 71986 39686 72038 39738
rect 72050 39686 72102 39738
rect 72114 39686 72166 39738
rect 63408 39584 63460 39636
rect 65524 39584 65576 39636
rect 66260 39584 66312 39636
rect 67548 39380 67600 39432
rect 74210 39142 74262 39194
rect 74274 39142 74326 39194
rect 74338 39142 74390 39194
rect 74402 39142 74454 39194
rect 74466 39142 74518 39194
rect 65248 39040 65300 39092
rect 63408 38884 63460 38936
rect 69848 38836 69900 38888
rect 65432 38700 65484 38752
rect 71858 38598 71910 38650
rect 71922 38598 71974 38650
rect 71986 38598 72038 38650
rect 72050 38598 72102 38650
rect 72114 38598 72166 38650
rect 69296 38496 69348 38548
rect 65984 38428 66036 38480
rect 66260 38428 66312 38480
rect 69480 38292 69532 38344
rect 74210 38054 74262 38106
rect 74274 38054 74326 38106
rect 74338 38054 74390 38106
rect 74402 38054 74454 38106
rect 74466 38054 74518 38106
rect 69112 37952 69164 38004
rect 70032 37748 70084 37800
rect 71858 37510 71910 37562
rect 71922 37510 71974 37562
rect 71986 37510 72038 37562
rect 72050 37510 72102 37562
rect 72114 37510 72166 37562
rect 65156 37340 65208 37392
rect 65616 37247 65668 37256
rect 65616 37213 65625 37247
rect 65625 37213 65659 37247
rect 65659 37213 65668 37247
rect 65616 37204 65668 37213
rect 67456 37204 67508 37256
rect 74210 36966 74262 37018
rect 74274 36966 74326 37018
rect 74338 36966 74390 37018
rect 74402 36966 74454 37018
rect 74466 36966 74518 37018
rect 65524 36864 65576 36916
rect 64972 36728 65024 36780
rect 65524 36728 65576 36780
rect 66904 36660 66956 36712
rect 64972 36524 65024 36576
rect 71858 36422 71910 36474
rect 71922 36422 71974 36474
rect 71986 36422 72038 36474
rect 72050 36422 72102 36474
rect 72114 36422 72166 36474
rect 64880 36320 64932 36372
rect 66352 36363 66404 36372
rect 66352 36329 66361 36363
rect 66361 36329 66395 36363
rect 66395 36329 66404 36363
rect 66352 36320 66404 36329
rect 67364 36184 67416 36236
rect 65984 36116 66036 36168
rect 68284 36116 68336 36168
rect 74210 35878 74262 35930
rect 74274 35878 74326 35930
rect 74338 35878 74390 35930
rect 74402 35878 74454 35930
rect 74466 35878 74518 35930
rect 66996 35776 67048 35828
rect 69388 35708 69440 35760
rect 64144 35640 64196 35692
rect 68376 35572 68428 35624
rect 71858 35334 71910 35386
rect 71922 35334 71974 35386
rect 71986 35334 72038 35386
rect 72050 35334 72102 35386
rect 72114 35334 72166 35386
rect 67916 35232 67968 35284
rect 64880 35164 64932 35216
rect 65156 35164 65208 35216
rect 69020 35096 69072 35148
rect 68468 35028 68520 35080
rect 65616 35003 65668 35012
rect 65616 34969 65625 35003
rect 65625 34969 65659 35003
rect 65659 34969 65668 35003
rect 65616 34960 65668 34969
rect 74210 34790 74262 34842
rect 74274 34790 74326 34842
rect 74338 34790 74390 34842
rect 74402 34790 74454 34842
rect 74466 34790 74518 34842
rect 65064 34688 65116 34740
rect 66812 34688 66864 34740
rect 67272 34620 67324 34672
rect 65064 34484 65116 34536
rect 66352 34484 66404 34536
rect 66812 34484 66864 34536
rect 67732 34527 67784 34536
rect 67732 34493 67741 34527
rect 67741 34493 67775 34527
rect 67775 34493 67784 34527
rect 67732 34484 67784 34493
rect 71858 34246 71910 34298
rect 71922 34246 71974 34298
rect 71986 34246 72038 34298
rect 72050 34246 72102 34298
rect 72114 34246 72166 34298
rect 65708 34144 65760 34196
rect 66260 34144 66312 34196
rect 67640 34144 67692 34196
rect 67088 34008 67140 34060
rect 65156 33940 65208 33992
rect 66996 33983 67048 33992
rect 66996 33949 67005 33983
rect 67005 33949 67039 33983
rect 67039 33949 67048 33983
rect 66996 33940 67048 33949
rect 68836 33940 68888 33992
rect 74210 33702 74262 33754
rect 74274 33702 74326 33754
rect 74338 33702 74390 33754
rect 74402 33702 74454 33754
rect 74466 33702 74518 33754
rect 65524 33600 65576 33652
rect 65708 33396 65760 33448
rect 64880 33260 64932 33312
rect 71858 33158 71910 33210
rect 71922 33158 71974 33210
rect 71986 33158 72038 33210
rect 72050 33158 72102 33210
rect 72114 33158 72166 33210
rect 66168 33056 66220 33108
rect 69296 32852 69348 32904
rect 74210 32614 74262 32666
rect 74274 32614 74326 32666
rect 74338 32614 74390 32666
rect 74402 32614 74454 32666
rect 74466 32614 74518 32666
rect 69572 32512 69624 32564
rect 70216 32308 70268 32360
rect 65248 32172 65300 32224
rect 71858 32070 71910 32122
rect 71922 32070 71974 32122
rect 71986 32070 72038 32122
rect 72050 32070 72102 32122
rect 72114 32070 72166 32122
rect 69664 31968 69716 32020
rect 67272 31900 67324 31952
rect 67824 31764 67876 31816
rect 74210 31526 74262 31578
rect 74274 31526 74326 31578
rect 74338 31526 74390 31578
rect 74402 31526 74454 31578
rect 74466 31526 74518 31578
rect 65340 31424 65392 31476
rect 69388 31220 69440 31272
rect 64880 31084 64932 31136
rect 71858 30982 71910 31034
rect 71922 30982 71974 31034
rect 71986 30982 72038 31034
rect 72050 30982 72102 31034
rect 72114 30982 72166 31034
rect 67180 30880 67232 30932
rect 69664 30676 69716 30728
rect 74210 30438 74262 30490
rect 74274 30438 74326 30490
rect 74338 30438 74390 30490
rect 74402 30438 74454 30490
rect 74466 30438 74518 30490
rect 65432 30268 65484 30320
rect 67180 30132 67232 30184
rect 65340 29996 65392 30048
rect 66260 29996 66312 30048
rect 66720 29996 66772 30048
rect 71858 29894 71910 29946
rect 71922 29894 71974 29946
rect 71986 29894 72038 29946
rect 72050 29894 72102 29946
rect 72114 29894 72166 29946
rect 66444 29792 66496 29844
rect 66168 29588 66220 29640
rect 66444 29520 66496 29572
rect 74210 29350 74262 29402
rect 74274 29350 74326 29402
rect 74338 29350 74390 29402
rect 74402 29350 74454 29402
rect 74466 29350 74518 29402
rect 66260 29291 66312 29300
rect 66260 29257 66269 29291
rect 66269 29257 66303 29291
rect 66303 29257 66312 29291
rect 66260 29248 66312 29257
rect 69572 29112 69624 29164
rect 66352 29044 66404 29096
rect 67272 29044 67324 29096
rect 65156 28976 65208 29028
rect 67272 28908 67324 28960
rect 71858 28806 71910 28858
rect 71922 28806 71974 28858
rect 71986 28806 72038 28858
rect 72050 28806 72102 28858
rect 72114 28806 72166 28858
rect 65616 28704 65668 28756
rect 69112 28704 69164 28756
rect 64880 28636 64932 28688
rect 66628 28432 66680 28484
rect 74210 28262 74262 28314
rect 74274 28262 74326 28314
rect 74338 28262 74390 28314
rect 74402 28262 74454 28314
rect 74466 28262 74518 28314
rect 65984 28160 66036 28212
rect 68008 27956 68060 28008
rect 65524 27820 65576 27872
rect 66628 27863 66680 27872
rect 66628 27829 66637 27863
rect 66637 27829 66671 27863
rect 66671 27829 66680 27863
rect 66628 27820 66680 27829
rect 69020 27820 69072 27872
rect 71858 27718 71910 27770
rect 71922 27718 71974 27770
rect 71986 27718 72038 27770
rect 72050 27718 72102 27770
rect 72114 27718 72166 27770
rect 65156 27616 65208 27668
rect 66720 27548 66772 27600
rect 64236 27480 64288 27532
rect 65800 27412 65852 27464
rect 69756 27344 69808 27396
rect 74210 27174 74262 27226
rect 74274 27174 74326 27226
rect 74338 27174 74390 27226
rect 74402 27174 74454 27226
rect 74466 27174 74518 27226
rect 67272 27072 67324 27124
rect 66536 27047 66588 27056
rect 66536 27013 66545 27047
rect 66545 27013 66579 27047
rect 66579 27013 66588 27047
rect 66536 27004 66588 27013
rect 64328 26936 64380 26988
rect 68744 26868 68796 26920
rect 64880 26732 64932 26784
rect 66444 26732 66496 26784
rect 71858 26630 71910 26682
rect 71922 26630 71974 26682
rect 71986 26630 72038 26682
rect 72050 26630 72102 26682
rect 72114 26630 72166 26682
rect 69204 26528 69256 26580
rect 67272 26324 67324 26376
rect 74210 26086 74262 26138
rect 74274 26086 74326 26138
rect 74338 26086 74390 26138
rect 74402 26086 74454 26138
rect 74466 26086 74518 26138
rect 69848 25984 69900 26036
rect 71504 25780 71556 25832
rect 65432 25644 65484 25696
rect 71858 25542 71910 25594
rect 71922 25542 71974 25594
rect 71986 25542 72038 25594
rect 72050 25542 72102 25594
rect 72114 25542 72166 25594
rect 67456 25440 67508 25492
rect 67088 25372 67140 25424
rect 67456 25304 67508 25356
rect 65984 25236 66036 25288
rect 67088 25236 67140 25288
rect 74210 24998 74262 25050
rect 74274 24998 74326 25050
rect 74338 24998 74390 25050
rect 74402 24998 74454 25050
rect 74466 24998 74518 25050
rect 65616 24828 65668 24880
rect 66260 24828 66312 24880
rect 66352 24803 66404 24812
rect 66352 24769 66361 24803
rect 66361 24769 66395 24803
rect 66395 24769 66404 24803
rect 66352 24760 66404 24769
rect 66260 24735 66312 24744
rect 66260 24701 66269 24735
rect 66269 24701 66303 24735
rect 66303 24701 66312 24735
rect 66260 24692 66312 24701
rect 69756 24692 69808 24744
rect 67364 24624 67416 24676
rect 71858 24454 71910 24506
rect 71922 24454 71974 24506
rect 71986 24454 72038 24506
rect 72050 24454 72102 24506
rect 72114 24454 72166 24506
rect 66904 24352 66956 24404
rect 68376 24352 68428 24404
rect 64880 24284 64932 24336
rect 66536 24216 66588 24268
rect 66352 24191 66404 24200
rect 66352 24157 66361 24191
rect 66361 24157 66395 24191
rect 66395 24157 66404 24191
rect 66352 24148 66404 24157
rect 74210 23910 74262 23962
rect 74274 23910 74326 23962
rect 74338 23910 74390 23962
rect 74402 23910 74454 23962
rect 74466 23910 74518 23962
rect 65616 23851 65668 23860
rect 65616 23817 65625 23851
rect 65625 23817 65659 23851
rect 65659 23817 65668 23851
rect 65616 23808 65668 23817
rect 66812 23808 66864 23860
rect 67732 23808 67784 23860
rect 64880 23672 64932 23724
rect 65616 23672 65668 23724
rect 66628 23604 66680 23656
rect 66812 23604 66864 23656
rect 68928 23604 68980 23656
rect 64880 23468 64932 23520
rect 71858 23366 71910 23418
rect 71922 23366 71974 23418
rect 71986 23366 72038 23418
rect 72050 23366 72102 23418
rect 72114 23366 72166 23418
rect 66720 23264 66772 23316
rect 66996 23196 67048 23248
rect 67364 23128 67416 23180
rect 66904 23103 66956 23112
rect 66904 23069 66913 23103
rect 66913 23069 66947 23103
rect 66947 23069 66956 23103
rect 66904 23060 66956 23069
rect 67916 23060 67968 23112
rect 65432 22992 65484 23044
rect 67456 22992 67508 23044
rect 74210 22822 74262 22874
rect 74274 22822 74326 22874
rect 74338 22822 74390 22874
rect 74402 22822 74454 22874
rect 74466 22822 74518 22874
rect 65708 22720 65760 22772
rect 66720 22516 66772 22568
rect 71858 22278 71910 22330
rect 71922 22278 71974 22330
rect 71986 22278 72038 22330
rect 72050 22278 72102 22330
rect 72114 22278 72166 22330
rect 65708 22108 65760 22160
rect 66444 22083 66496 22092
rect 66444 22049 66453 22083
rect 66453 22049 66487 22083
rect 66487 22049 66496 22083
rect 66444 22040 66496 22049
rect 68560 22040 68612 22092
rect 70124 22083 70176 22092
rect 70124 22049 70133 22083
rect 70133 22049 70167 22083
rect 70167 22049 70176 22083
rect 70124 22040 70176 22049
rect 67640 21972 67692 22024
rect 69940 21972 69992 22024
rect 71596 21972 71648 22024
rect 74210 21734 74262 21786
rect 74274 21734 74326 21786
rect 74338 21734 74390 21786
rect 74402 21734 74454 21786
rect 74466 21734 74518 21786
rect 65156 21632 65208 21684
rect 69848 21428 69900 21480
rect 65156 21360 65208 21412
rect 65524 21360 65576 21412
rect 64788 21292 64840 21344
rect 71858 21190 71910 21242
rect 71922 21190 71974 21242
rect 71986 21190 72038 21242
rect 72050 21190 72102 21242
rect 72114 21190 72166 21242
rect 68192 21131 68244 21140
rect 68192 21097 68201 21131
rect 68201 21097 68235 21131
rect 68235 21097 68244 21131
rect 68192 21088 68244 21097
rect 65616 20884 65668 20936
rect 70124 20884 70176 20936
rect 66260 20748 66312 20800
rect 67456 20748 67508 20800
rect 74210 20646 74262 20698
rect 74274 20646 74326 20698
rect 74338 20646 74390 20698
rect 74402 20646 74454 20698
rect 74466 20646 74518 20698
rect 67548 20544 67600 20596
rect 69480 20476 69532 20528
rect 68284 20408 68336 20460
rect 68376 20340 68428 20392
rect 65708 20272 65760 20324
rect 66996 20272 67048 20324
rect 70032 20204 70084 20256
rect 71858 20102 71910 20154
rect 71922 20102 71974 20154
rect 71986 20102 72038 20154
rect 72050 20102 72102 20154
rect 72114 20102 72166 20154
rect 65984 20000 66036 20052
rect 66628 19932 66680 19984
rect 67088 19932 67140 19984
rect 65524 19864 65576 19916
rect 65984 19864 66036 19916
rect 69480 19796 69532 19848
rect 74210 19558 74262 19610
rect 74274 19558 74326 19610
rect 74338 19558 74390 19610
rect 74402 19558 74454 19610
rect 74466 19558 74518 19610
rect 68192 19456 68244 19508
rect 68560 19252 68612 19304
rect 72332 19184 72384 19236
rect 71858 19014 71910 19066
rect 71922 19014 71974 19066
rect 71986 19014 72038 19066
rect 72050 19014 72102 19066
rect 72114 19014 72166 19066
rect 68468 18912 68520 18964
rect 65524 18708 65576 18760
rect 72424 18708 72476 18760
rect 74210 18470 74262 18522
rect 74274 18470 74326 18522
rect 74338 18470 74390 18522
rect 74402 18470 74454 18522
rect 74466 18470 74518 18522
rect 65432 18368 65484 18420
rect 64880 18232 64932 18284
rect 65432 18232 65484 18284
rect 69204 18164 69256 18216
rect 65708 18028 65760 18080
rect 71858 17926 71910 17978
rect 71922 17926 71974 17978
rect 71986 17926 72038 17978
rect 72050 17926 72102 17978
rect 72114 17926 72166 17978
rect 68836 17824 68888 17876
rect 70584 17620 70636 17672
rect 74210 17382 74262 17434
rect 74274 17382 74326 17434
rect 74338 17382 74390 17434
rect 74402 17382 74454 17434
rect 74466 17382 74518 17434
rect 65616 17323 65668 17332
rect 65616 17289 65625 17323
rect 65625 17289 65659 17323
rect 65659 17289 65668 17323
rect 65616 17280 65668 17289
rect 70216 17280 70268 17332
rect 70492 17144 70544 17196
rect 66260 17119 66312 17128
rect 66260 17085 66269 17119
rect 66269 17085 66303 17119
rect 66303 17085 66312 17119
rect 66260 17076 66312 17085
rect 72240 17076 72292 17128
rect 71858 16838 71910 16890
rect 71922 16838 71974 16890
rect 71986 16838 72038 16890
rect 72050 16838 72102 16890
rect 72114 16838 72166 16890
rect 64880 16600 64932 16652
rect 72516 16600 72568 16652
rect 67824 16532 67876 16584
rect 74210 16294 74262 16346
rect 74274 16294 74326 16346
rect 74338 16294 74390 16346
rect 74402 16294 74454 16346
rect 74466 16294 74518 16346
rect 66168 16192 66220 16244
rect 64696 16056 64748 16108
rect 66996 16056 67048 16108
rect 70400 15988 70452 16040
rect 71858 15750 71910 15802
rect 71922 15750 71974 15802
rect 71986 15750 72038 15802
rect 72050 15750 72102 15802
rect 72114 15750 72166 15802
rect 69664 15648 69716 15700
rect 65616 15512 65668 15564
rect 70952 15444 71004 15496
rect 65708 15308 65760 15360
rect 66260 15308 66312 15360
rect 67548 15308 67600 15360
rect 70768 15308 70820 15360
rect 74210 15206 74262 15258
rect 74274 15206 74326 15258
rect 74338 15206 74390 15258
rect 74402 15206 74454 15258
rect 74466 15206 74518 15258
rect 69572 15104 69624 15156
rect 69664 14900 69716 14952
rect 72608 14832 72660 14884
rect 71858 14662 71910 14714
rect 71922 14662 71974 14714
rect 71986 14662 72038 14714
rect 72050 14662 72102 14714
rect 72114 14662 72166 14714
rect 65524 14560 65576 14612
rect 69388 14492 69440 14544
rect 69572 14492 69624 14544
rect 65616 14356 65668 14408
rect 67732 14356 67784 14408
rect 74210 14118 74262 14170
rect 74274 14118 74326 14170
rect 74338 14118 74390 14170
rect 74402 14118 74454 14170
rect 74466 14118 74518 14170
rect 71858 13574 71910 13626
rect 71922 13574 71974 13626
rect 71986 13574 72038 13626
rect 72050 13574 72102 13626
rect 72114 13574 72166 13626
rect 64880 13472 64932 13524
rect 64880 13336 64932 13388
rect 65524 13336 65576 13388
rect 68100 13268 68152 13320
rect 74210 13030 74262 13082
rect 74274 13030 74326 13082
rect 74338 13030 74390 13082
rect 74402 13030 74454 13082
rect 74466 13030 74518 13082
rect 65524 12724 65576 12776
rect 66168 12588 66220 12640
rect 71858 12486 71910 12538
rect 71922 12486 71974 12538
rect 71986 12486 72038 12538
rect 72050 12486 72102 12538
rect 72114 12486 72166 12538
rect 74210 11942 74262 11994
rect 74274 11942 74326 11994
rect 74338 11942 74390 11994
rect 74402 11942 74454 11994
rect 74466 11942 74518 11994
rect 65616 11883 65668 11892
rect 65616 11849 65625 11883
rect 65625 11849 65659 11883
rect 65659 11849 65668 11883
rect 65616 11840 65668 11849
rect 69204 11636 69256 11688
rect 64972 11500 65024 11552
rect 65524 11500 65576 11552
rect 63868 11432 63920 11484
rect 64512 11432 64564 11484
rect 63500 11364 63552 11416
rect 64328 11364 64380 11416
rect 71858 11398 71910 11450
rect 71922 11398 71974 11450
rect 71986 11398 72038 11450
rect 72050 11398 72102 11450
rect 72114 11398 72166 11450
rect 63592 11296 63644 11348
rect 63868 11296 63920 11348
rect 64972 11228 65024 11280
rect 63408 11092 63460 11144
rect 70860 11092 70912 11144
rect 74210 10854 74262 10906
rect 74274 10854 74326 10906
rect 74338 10854 74390 10906
rect 74402 10854 74454 10906
rect 74466 10854 74518 10906
rect 64880 10548 64932 10600
rect 65616 10548 65668 10600
rect 65616 10412 65668 10464
rect 63500 10292 63552 10344
rect 71858 10310 71910 10362
rect 71922 10310 71974 10362
rect 71986 10310 72038 10362
rect 72050 10310 72102 10362
rect 72114 10310 72166 10362
rect 74210 9766 74262 9818
rect 74274 9766 74326 9818
rect 74338 9766 74390 9818
rect 74402 9766 74454 9818
rect 74466 9766 74518 9818
rect 64972 9324 65024 9376
rect 71858 9222 71910 9274
rect 71922 9222 71974 9274
rect 71986 9222 72038 9274
rect 72050 9222 72102 9274
rect 72114 9222 72166 9274
rect 74210 8678 74262 8730
rect 74274 8678 74326 8730
rect 74338 8678 74390 8730
rect 74402 8678 74454 8730
rect 74466 8678 74518 8730
rect 71858 8134 71910 8186
rect 71922 8134 71974 8186
rect 71986 8134 72038 8186
rect 72050 8134 72102 8186
rect 72114 8134 72166 8186
rect 59184 7828 59236 7880
rect 67548 8032 67600 8084
rect 63224 7828 63276 7880
rect 66812 7964 66864 8016
rect 64880 7828 64932 7880
rect 65156 7828 65208 7880
rect 47308 7760 47360 7812
rect 55772 7760 55824 7812
rect 59560 7760 59612 7812
rect 63408 7760 63460 7812
rect 44824 7692 44876 7744
rect 66352 7760 66404 7812
rect 65156 7692 65208 7744
rect 65340 7692 65392 7744
rect 33048 7556 33100 7608
rect 63592 7556 63644 7608
rect 74210 7590 74262 7642
rect 74274 7590 74326 7642
rect 74338 7590 74390 7642
rect 74402 7590 74454 7642
rect 74466 7590 74518 7642
rect 55772 7420 55824 7472
rect 67180 7488 67232 7540
rect 63132 7420 63184 7472
rect 65800 7420 65852 7472
rect 62672 7352 62724 7404
rect 67456 7352 67508 7404
rect 62304 7284 62356 7336
rect 66076 7284 66128 7336
rect 55036 7216 55088 7268
rect 64236 7216 64288 7268
rect 62764 7148 62816 7200
rect 68744 7148 68796 7200
rect 58624 7012 58676 7064
rect 64512 7012 64564 7064
rect 71858 7046 71910 7098
rect 71922 7046 71974 7098
rect 71986 7046 72038 7098
rect 72050 7046 72102 7098
rect 72114 7046 72166 7098
rect 63316 6944 63368 6996
rect 67916 6944 67968 6996
rect 61476 6876 61528 6928
rect 63500 6876 63552 6928
rect 49056 6808 49108 6860
rect 49792 6740 49844 6792
rect 55772 6740 55824 6792
rect 56508 6808 56560 6860
rect 70400 6808 70452 6860
rect 66904 6740 66956 6792
rect 47768 6604 47820 6656
rect 66720 6672 66772 6724
rect 55956 6604 56008 6656
rect 60924 6604 60976 6656
rect 61108 6604 61160 6656
rect 68928 6604 68980 6656
rect 49608 6536 49660 6588
rect 62764 6536 62816 6588
rect 36728 6468 36780 6520
rect 63132 6468 63184 6520
rect 74210 6502 74262 6554
rect 74274 6502 74326 6554
rect 74338 6502 74390 6554
rect 74402 6502 74454 6554
rect 74466 6502 74518 6554
rect 48228 6400 48280 6452
rect 46756 6332 46808 6384
rect 61108 6332 61160 6384
rect 68008 6400 68060 6452
rect 42248 6264 42300 6316
rect 65800 6332 65852 6384
rect 69848 6332 69900 6384
rect 67364 6264 67416 6316
rect 50712 6196 50764 6248
rect 63316 6196 63368 6248
rect 63592 6196 63644 6248
rect 64328 6196 64380 6248
rect 56324 6128 56376 6180
rect 64972 6128 65024 6180
rect 56232 6060 56284 6112
rect 69204 6060 69256 6112
rect 71858 5958 71910 6010
rect 71922 5958 71974 6010
rect 71986 5958 72038 6010
rect 72050 5958 72102 6010
rect 72114 5958 72166 6010
rect 39488 5899 39540 5908
rect 39488 5865 39497 5899
rect 39497 5865 39531 5899
rect 39531 5865 39540 5899
rect 39488 5856 39540 5865
rect 41696 5899 41748 5908
rect 41696 5865 41705 5899
rect 41705 5865 41739 5899
rect 41739 5865 41748 5899
rect 41696 5856 41748 5865
rect 49608 5899 49660 5908
rect 49608 5865 49617 5899
rect 49617 5865 49651 5899
rect 49651 5865 49660 5899
rect 49608 5856 49660 5865
rect 50712 5899 50764 5908
rect 50712 5865 50721 5899
rect 50721 5865 50755 5899
rect 50755 5865 50764 5899
rect 50712 5856 50764 5865
rect 40408 5831 40460 5840
rect 40408 5797 40417 5831
rect 40417 5797 40451 5831
rect 40451 5797 40460 5831
rect 40408 5788 40460 5797
rect 41604 5788 41656 5840
rect 61108 5856 61160 5908
rect 72240 5856 72292 5908
rect 32312 5720 32364 5772
rect 44732 5720 44784 5772
rect 28908 5695 28960 5704
rect 28908 5661 28917 5695
rect 28917 5661 28951 5695
rect 28951 5661 28960 5695
rect 28908 5652 28960 5661
rect 29552 5652 29604 5704
rect 30380 5652 30432 5704
rect 30748 5652 30800 5704
rect 31392 5695 31444 5704
rect 31392 5661 31401 5695
rect 31401 5661 31435 5695
rect 31435 5661 31444 5695
rect 31392 5652 31444 5661
rect 35164 5652 35216 5704
rect 36452 5695 36504 5704
rect 36452 5661 36461 5695
rect 36461 5661 36495 5695
rect 36495 5661 36504 5695
rect 36452 5652 36504 5661
rect 36728 5695 36780 5704
rect 36728 5661 36737 5695
rect 36737 5661 36771 5695
rect 36771 5661 36780 5695
rect 36728 5652 36780 5661
rect 37188 5695 37240 5704
rect 37188 5661 37197 5695
rect 37197 5661 37231 5695
rect 37231 5661 37240 5695
rect 37188 5652 37240 5661
rect 38108 5695 38160 5704
rect 38108 5661 38117 5695
rect 38117 5661 38151 5695
rect 38151 5661 38160 5695
rect 38108 5652 38160 5661
rect 38752 5695 38804 5704
rect 38752 5661 38761 5695
rect 38761 5661 38795 5695
rect 38795 5661 38804 5695
rect 38752 5652 38804 5661
rect 38844 5695 38896 5704
rect 38844 5661 38853 5695
rect 38853 5661 38887 5695
rect 38887 5661 38896 5695
rect 38844 5652 38896 5661
rect 39764 5695 39816 5704
rect 39764 5661 39773 5695
rect 39773 5661 39807 5695
rect 39807 5661 39816 5695
rect 39764 5652 39816 5661
rect 40408 5652 40460 5704
rect 42708 5652 42760 5704
rect 29368 5516 29420 5568
rect 30840 5559 30892 5568
rect 30840 5525 30849 5559
rect 30849 5525 30883 5559
rect 30883 5525 30892 5559
rect 30840 5516 30892 5525
rect 38936 5584 38988 5636
rect 48964 5695 49016 5704
rect 48964 5661 48973 5695
rect 48973 5661 49007 5695
rect 49007 5661 49016 5695
rect 48964 5652 49016 5661
rect 49700 5652 49752 5704
rect 50804 5695 50856 5704
rect 50804 5661 50813 5695
rect 50813 5661 50847 5695
rect 50847 5661 50856 5695
rect 50804 5652 50856 5661
rect 51540 5695 51592 5704
rect 51540 5661 51549 5695
rect 51549 5661 51583 5695
rect 51583 5661 51592 5695
rect 51540 5652 51592 5661
rect 52460 5652 52512 5704
rect 53840 5652 53892 5704
rect 55036 5695 55088 5704
rect 55036 5661 55045 5695
rect 55045 5661 55079 5695
rect 55079 5661 55088 5695
rect 55036 5652 55088 5661
rect 56324 5695 56376 5704
rect 56324 5661 56333 5695
rect 56333 5661 56367 5695
rect 56367 5661 56376 5695
rect 56324 5652 56376 5661
rect 56692 5695 56744 5704
rect 56692 5661 56701 5695
rect 56701 5661 56735 5695
rect 56735 5661 56744 5695
rect 56692 5652 56744 5661
rect 60280 5720 60332 5772
rect 60464 5763 60516 5772
rect 60464 5729 60473 5763
rect 60473 5729 60507 5763
rect 60507 5729 60516 5763
rect 60464 5720 60516 5729
rect 71504 5788 71556 5840
rect 61292 5720 61344 5772
rect 61384 5720 61436 5772
rect 69756 5720 69808 5772
rect 67640 5652 67692 5704
rect 60280 5584 60332 5636
rect 69480 5584 69532 5636
rect 37280 5516 37332 5568
rect 45468 5516 45520 5568
rect 58532 5516 58584 5568
rect 66168 5516 66220 5568
rect 69940 5516 69992 5568
rect 71136 5516 71188 5568
rect 71596 5516 71648 5568
rect 73436 5516 73488 5568
rect 4210 5414 4262 5466
rect 4274 5414 4326 5466
rect 4338 5414 4390 5466
rect 4402 5414 4454 5466
rect 4466 5414 4518 5466
rect 14210 5414 14262 5466
rect 14274 5414 14326 5466
rect 14338 5414 14390 5466
rect 14402 5414 14454 5466
rect 14466 5414 14518 5466
rect 24210 5414 24262 5466
rect 24274 5414 24326 5466
rect 24338 5414 24390 5466
rect 24402 5414 24454 5466
rect 24466 5414 24518 5466
rect 34210 5414 34262 5466
rect 34274 5414 34326 5466
rect 34338 5414 34390 5466
rect 34402 5414 34454 5466
rect 34466 5414 34518 5466
rect 44210 5414 44262 5466
rect 44274 5414 44326 5466
rect 44338 5414 44390 5466
rect 44402 5414 44454 5466
rect 44466 5414 44518 5466
rect 54210 5414 54262 5466
rect 54274 5414 54326 5466
rect 54338 5414 54390 5466
rect 54402 5414 54454 5466
rect 54466 5414 54518 5466
rect 64210 5414 64262 5466
rect 64274 5414 64326 5466
rect 64338 5414 64390 5466
rect 64402 5414 64454 5466
rect 64466 5414 64518 5466
rect 74210 5414 74262 5466
rect 74274 5414 74326 5466
rect 74338 5414 74390 5466
rect 74402 5414 74454 5466
rect 74466 5414 74518 5466
rect 36452 5312 36504 5364
rect 41604 5312 41656 5364
rect 42708 5312 42760 5364
rect 42892 5312 42944 5364
rect 38108 5244 38160 5296
rect 42248 5244 42300 5296
rect 46112 5287 46164 5296
rect 46112 5253 46121 5287
rect 46121 5253 46155 5287
rect 46155 5253 46164 5287
rect 46112 5244 46164 5253
rect 47308 5355 47360 5364
rect 47308 5321 47317 5355
rect 47317 5321 47351 5355
rect 47351 5321 47360 5355
rect 47308 5312 47360 5321
rect 48228 5355 48280 5364
rect 48228 5321 48237 5355
rect 48237 5321 48271 5355
rect 48271 5321 48280 5355
rect 48228 5312 48280 5321
rect 49056 5355 49108 5364
rect 49056 5321 49065 5355
rect 49065 5321 49099 5355
rect 49099 5321 49108 5355
rect 49056 5312 49108 5321
rect 49792 5355 49844 5364
rect 49792 5321 49801 5355
rect 49801 5321 49835 5355
rect 49835 5321 49844 5355
rect 49792 5312 49844 5321
rect 53472 5312 53524 5364
rect 54024 5355 54076 5364
rect 54024 5321 54033 5355
rect 54033 5321 54067 5355
rect 54067 5321 54076 5355
rect 54024 5312 54076 5321
rect 48964 5244 49016 5296
rect 29184 5219 29236 5228
rect 29184 5185 29193 5219
rect 29193 5185 29227 5219
rect 29227 5185 29236 5219
rect 29184 5176 29236 5185
rect 29368 5219 29420 5228
rect 29368 5185 29377 5219
rect 29377 5185 29411 5219
rect 29411 5185 29420 5219
rect 29368 5176 29420 5185
rect 32220 5176 32272 5228
rect 37280 5176 37332 5228
rect 25044 5108 25096 5160
rect 26148 5108 26200 5160
rect 28356 5108 28408 5160
rect 31300 5108 31352 5160
rect 33416 5151 33468 5160
rect 33416 5117 33425 5151
rect 33425 5117 33459 5151
rect 33459 5117 33468 5151
rect 33416 5108 33468 5117
rect 33784 5108 33836 5160
rect 36544 5108 36596 5160
rect 37740 5108 37792 5160
rect 44088 5219 44140 5228
rect 44088 5185 44097 5219
rect 44097 5185 44131 5219
rect 44131 5185 44140 5219
rect 44088 5176 44140 5185
rect 44732 5219 44784 5228
rect 44732 5185 44741 5219
rect 44741 5185 44775 5219
rect 44775 5185 44784 5219
rect 44732 5176 44784 5185
rect 45468 5219 45520 5228
rect 45468 5185 45477 5219
rect 45477 5185 45511 5219
rect 45511 5185 45520 5219
rect 45468 5176 45520 5185
rect 46204 5176 46256 5228
rect 52828 5176 52880 5228
rect 55864 5244 55916 5296
rect 60372 5312 60424 5364
rect 67732 5312 67784 5364
rect 60556 5244 60608 5296
rect 69296 5244 69348 5296
rect 56600 5176 56652 5228
rect 69112 5176 69164 5228
rect 39212 5151 39264 5160
rect 39212 5117 39221 5151
rect 39221 5117 39255 5151
rect 39255 5117 39264 5151
rect 39212 5108 39264 5117
rect 40132 5151 40184 5160
rect 40132 5117 40141 5151
rect 40141 5117 40175 5151
rect 40175 5117 40184 5151
rect 40132 5108 40184 5117
rect 46664 5151 46716 5160
rect 46664 5117 46673 5151
rect 46673 5117 46707 5151
rect 46707 5117 46716 5151
rect 46664 5108 46716 5117
rect 47584 5151 47636 5160
rect 47584 5117 47593 5151
rect 47593 5117 47627 5151
rect 47627 5117 47636 5151
rect 47584 5108 47636 5117
rect 48412 5151 48464 5160
rect 48412 5117 48421 5151
rect 48421 5117 48455 5151
rect 48455 5117 48464 5151
rect 48412 5108 48464 5117
rect 49148 5151 49200 5160
rect 49148 5117 49157 5151
rect 49157 5117 49191 5151
rect 49191 5117 49200 5151
rect 49148 5108 49200 5117
rect 49792 5108 49844 5160
rect 50160 5108 50212 5160
rect 51264 5151 51316 5160
rect 51264 5117 51273 5151
rect 51273 5117 51307 5151
rect 51307 5117 51316 5151
rect 51264 5108 51316 5117
rect 51356 5151 51408 5160
rect 51356 5117 51365 5151
rect 51365 5117 51399 5151
rect 51399 5117 51408 5151
rect 51356 5108 51408 5117
rect 51724 5108 51776 5160
rect 53288 5151 53340 5160
rect 53288 5117 53297 5151
rect 53297 5117 53331 5151
rect 53331 5117 53340 5151
rect 53288 5108 53340 5117
rect 53380 5151 53432 5160
rect 53380 5117 53389 5151
rect 53389 5117 53423 5151
rect 53423 5117 53432 5151
rect 53380 5108 53432 5117
rect 53472 5108 53524 5160
rect 54852 5151 54904 5160
rect 54852 5117 54861 5151
rect 54861 5117 54895 5151
rect 54895 5117 54904 5151
rect 54852 5108 54904 5117
rect 55404 5108 55456 5160
rect 69572 5108 69624 5160
rect 23572 5040 23624 5092
rect 39948 5040 40000 5092
rect 43628 5040 43680 5092
rect 26700 5015 26752 5024
rect 26700 4981 26709 5015
rect 26709 4981 26743 5015
rect 26743 4981 26752 5015
rect 26700 4972 26752 4981
rect 27896 5015 27948 5024
rect 27896 4981 27905 5015
rect 27905 4981 27939 5015
rect 27939 4981 27948 5015
rect 27896 4972 27948 4981
rect 30656 5015 30708 5024
rect 30656 4981 30665 5015
rect 30665 4981 30699 5015
rect 30699 4981 30708 5015
rect 30656 4972 30708 4981
rect 31576 4972 31628 5024
rect 32864 5015 32916 5024
rect 32864 4981 32873 5015
rect 32873 4981 32907 5015
rect 32907 4981 32916 5015
rect 32864 4972 32916 4981
rect 36084 4972 36136 5024
rect 38844 4972 38896 5024
rect 69388 5040 69440 5092
rect 55496 5015 55548 5024
rect 55496 4981 55505 5015
rect 55505 4981 55539 5015
rect 55539 4981 55548 5015
rect 55496 4972 55548 4981
rect 56232 5015 56284 5024
rect 56232 4981 56241 5015
rect 56241 4981 56275 5015
rect 56275 4981 56284 5015
rect 56232 4972 56284 4981
rect 56416 4972 56468 5024
rect 63224 4972 63276 5024
rect 1858 4870 1910 4922
rect 1922 4870 1974 4922
rect 1986 4870 2038 4922
rect 2050 4870 2102 4922
rect 2114 4870 2166 4922
rect 11858 4870 11910 4922
rect 11922 4870 11974 4922
rect 11986 4870 12038 4922
rect 12050 4870 12102 4922
rect 12114 4870 12166 4922
rect 21858 4870 21910 4922
rect 21922 4870 21974 4922
rect 21986 4870 22038 4922
rect 22050 4870 22102 4922
rect 22114 4870 22166 4922
rect 31858 4870 31910 4922
rect 31922 4870 31974 4922
rect 31986 4870 32038 4922
rect 32050 4870 32102 4922
rect 32114 4870 32166 4922
rect 41858 4870 41910 4922
rect 41922 4870 41974 4922
rect 41986 4870 42038 4922
rect 42050 4870 42102 4922
rect 42114 4870 42166 4922
rect 51858 4870 51910 4922
rect 51922 4870 51974 4922
rect 51986 4870 52038 4922
rect 52050 4870 52102 4922
rect 52114 4870 52166 4922
rect 61858 4870 61910 4922
rect 61922 4870 61974 4922
rect 61986 4870 62038 4922
rect 62050 4870 62102 4922
rect 62114 4870 62166 4922
rect 71858 4870 71910 4922
rect 71922 4870 71974 4922
rect 71986 4870 72038 4922
rect 72050 4870 72102 4922
rect 72114 4870 72166 4922
rect 26148 4811 26200 4820
rect 26148 4777 26157 4811
rect 26157 4777 26191 4811
rect 26191 4777 26200 4811
rect 26148 4768 26200 4777
rect 31300 4811 31352 4820
rect 31300 4777 31309 4811
rect 31309 4777 31343 4811
rect 31343 4777 31352 4811
rect 31300 4768 31352 4777
rect 33784 4811 33836 4820
rect 33784 4777 33793 4811
rect 33793 4777 33827 4811
rect 33827 4777 33836 4811
rect 33784 4768 33836 4777
rect 29552 4700 29604 4752
rect 26332 4632 26384 4684
rect 24860 4564 24912 4616
rect 26240 4607 26292 4616
rect 26240 4573 26249 4607
rect 26249 4573 26283 4607
rect 26283 4573 26292 4607
rect 26240 4564 26292 4573
rect 28080 4564 28132 4616
rect 28632 4607 28684 4616
rect 28632 4573 28641 4607
rect 28641 4573 28675 4607
rect 28675 4573 28684 4607
rect 28632 4564 28684 4573
rect 29828 4607 29880 4616
rect 29828 4573 29837 4607
rect 29837 4573 29871 4607
rect 29871 4573 29880 4607
rect 29828 4564 29880 4573
rect 31300 4564 31352 4616
rect 29644 4496 29696 4548
rect 30932 4496 30984 4548
rect 32680 4564 32732 4616
rect 33140 4607 33192 4616
rect 33140 4573 33149 4607
rect 33149 4573 33183 4607
rect 33183 4573 33192 4607
rect 33140 4564 33192 4573
rect 33968 4607 34020 4616
rect 33968 4573 33977 4607
rect 33977 4573 34011 4607
rect 34011 4573 34020 4607
rect 33968 4564 34020 4573
rect 36084 4632 36136 4684
rect 40592 4743 40644 4752
rect 40592 4709 40601 4743
rect 40601 4709 40635 4743
rect 40635 4709 40644 4743
rect 40592 4700 40644 4709
rect 34612 4607 34664 4616
rect 34612 4573 34621 4607
rect 34621 4573 34655 4607
rect 34655 4573 34664 4607
rect 34612 4564 34664 4573
rect 35256 4539 35308 4548
rect 35256 4505 35265 4539
rect 35265 4505 35299 4539
rect 35299 4505 35308 4539
rect 35256 4496 35308 4505
rect 36360 4607 36412 4616
rect 36360 4573 36369 4607
rect 36369 4573 36403 4607
rect 36403 4573 36412 4607
rect 36360 4564 36412 4573
rect 37740 4564 37792 4616
rect 36912 4496 36964 4548
rect 38016 4539 38068 4548
rect 38016 4505 38025 4539
rect 38025 4505 38059 4539
rect 38059 4505 38068 4539
rect 38016 4496 38068 4505
rect 39948 4607 40000 4616
rect 39948 4573 39957 4607
rect 39957 4573 39991 4607
rect 39991 4573 40000 4607
rect 39948 4564 40000 4573
rect 40224 4564 40276 4616
rect 49148 4768 49200 4820
rect 54024 4768 54076 4820
rect 65708 4768 65760 4820
rect 43628 4700 43680 4752
rect 66444 4700 66496 4752
rect 67272 4632 67324 4684
rect 44088 4607 44140 4616
rect 44088 4573 44097 4607
rect 44097 4573 44131 4607
rect 44131 4573 44140 4607
rect 44088 4564 44140 4573
rect 44824 4564 44876 4616
rect 45008 4607 45060 4616
rect 45008 4573 45017 4607
rect 45017 4573 45051 4607
rect 45051 4573 45060 4607
rect 45008 4564 45060 4573
rect 45100 4564 45152 4616
rect 46756 4607 46808 4616
rect 46756 4573 46765 4607
rect 46765 4573 46799 4607
rect 46799 4573 46808 4607
rect 46756 4564 46808 4573
rect 47216 4607 47268 4616
rect 47216 4573 47225 4607
rect 47225 4573 47259 4607
rect 47259 4573 47268 4607
rect 47216 4564 47268 4573
rect 47768 4607 47820 4616
rect 47768 4573 47777 4607
rect 47777 4573 47811 4607
rect 47811 4573 47820 4607
rect 47768 4564 47820 4573
rect 47860 4607 47912 4616
rect 47860 4573 47869 4607
rect 47869 4573 47903 4607
rect 47903 4573 47912 4607
rect 47860 4564 47912 4573
rect 49608 4564 49660 4616
rect 53288 4564 53340 4616
rect 60556 4564 60608 4616
rect 66536 4496 66588 4548
rect 23480 4428 23532 4480
rect 27344 4471 27396 4480
rect 27344 4437 27353 4471
rect 27353 4437 27387 4471
rect 27387 4437 27396 4471
rect 27344 4428 27396 4437
rect 29276 4471 29328 4480
rect 29276 4437 29285 4471
rect 29285 4437 29319 4471
rect 29319 4437 29328 4471
rect 29276 4428 29328 4437
rect 30472 4471 30524 4480
rect 30472 4437 30481 4471
rect 30481 4437 30515 4471
rect 30515 4437 30524 4471
rect 30472 4428 30524 4437
rect 30564 4471 30616 4480
rect 30564 4437 30573 4471
rect 30573 4437 30607 4471
rect 30607 4437 30616 4471
rect 30564 4428 30616 4437
rect 32404 4471 32456 4480
rect 32404 4437 32413 4471
rect 32413 4437 32447 4471
rect 32447 4437 32456 4471
rect 32404 4428 32456 4437
rect 36728 4471 36780 4480
rect 36728 4437 36737 4471
rect 36737 4437 36771 4471
rect 36771 4437 36780 4471
rect 36728 4428 36780 4437
rect 37924 4471 37976 4480
rect 37924 4437 37933 4471
rect 37933 4437 37967 4471
rect 37967 4437 37976 4471
rect 37924 4428 37976 4437
rect 42892 4428 42944 4480
rect 45652 4471 45704 4480
rect 45652 4437 45661 4471
rect 45661 4437 45695 4471
rect 45695 4437 45704 4471
rect 45652 4428 45704 4437
rect 51724 4428 51776 4480
rect 56692 4428 56744 4480
rect 4210 4326 4262 4378
rect 4274 4326 4326 4378
rect 4338 4326 4390 4378
rect 4402 4326 4454 4378
rect 4466 4326 4518 4378
rect 14210 4326 14262 4378
rect 14274 4326 14326 4378
rect 14338 4326 14390 4378
rect 14402 4326 14454 4378
rect 14466 4326 14518 4378
rect 24210 4326 24262 4378
rect 24274 4326 24326 4378
rect 24338 4326 24390 4378
rect 24402 4326 24454 4378
rect 24466 4326 24518 4378
rect 34210 4326 34262 4378
rect 34274 4326 34326 4378
rect 34338 4326 34390 4378
rect 34402 4326 34454 4378
rect 34466 4326 34518 4378
rect 44210 4326 44262 4378
rect 44274 4326 44326 4378
rect 44338 4326 44390 4378
rect 44402 4326 44454 4378
rect 44466 4326 44518 4378
rect 54210 4326 54262 4378
rect 54274 4326 54326 4378
rect 54338 4326 54390 4378
rect 54402 4326 54454 4378
rect 54466 4326 54518 4378
rect 64210 4326 64262 4378
rect 64274 4326 64326 4378
rect 64338 4326 64390 4378
rect 64402 4326 64454 4378
rect 64466 4326 64518 4378
rect 74210 4326 74262 4378
rect 74274 4326 74326 4378
rect 74338 4326 74390 4378
rect 74402 4326 74454 4378
rect 74466 4326 74518 4378
rect 36728 4224 36780 4276
rect 43536 4224 43588 4276
rect 45652 4224 45704 4276
rect 56416 4224 56468 4276
rect 60464 4224 60516 4276
rect 63868 4224 63920 4276
rect 31116 4156 31168 4208
rect 32864 4156 32916 4208
rect 37924 4156 37976 4208
rect 26516 4088 26568 4140
rect 24584 4063 24636 4072
rect 24584 4029 24593 4063
rect 24593 4029 24627 4063
rect 24627 4029 24636 4063
rect 24584 4020 24636 4029
rect 25136 4020 25188 4072
rect 25964 4020 26016 4072
rect 27712 4020 27764 4072
rect 29184 4088 29236 4140
rect 29276 4088 29328 4140
rect 29644 4131 29696 4140
rect 29644 4097 29653 4131
rect 29653 4097 29687 4131
rect 29687 4097 29696 4131
rect 29644 4088 29696 4097
rect 30472 4088 30524 4140
rect 30656 4088 30708 4140
rect 32312 4088 32364 4140
rect 33140 4088 33192 4140
rect 33324 4088 33376 4140
rect 29368 4020 29420 4072
rect 30380 4063 30432 4072
rect 30380 4029 30389 4063
rect 30389 4029 30423 4063
rect 30423 4029 30432 4063
rect 30380 4020 30432 4029
rect 31024 4020 31076 4072
rect 32496 4020 32548 4072
rect 33876 4020 33928 4072
rect 34796 4020 34848 4072
rect 34980 4020 35032 4072
rect 35992 4063 36044 4072
rect 35992 4029 36001 4063
rect 36001 4029 36035 4063
rect 36035 4029 36044 4063
rect 35992 4020 36044 4029
rect 37832 4131 37884 4140
rect 37832 4097 37841 4131
rect 37841 4097 37875 4131
rect 37875 4097 37884 4131
rect 37832 4088 37884 4097
rect 38936 4131 38988 4140
rect 38936 4097 38945 4131
rect 38945 4097 38979 4131
rect 38979 4097 38988 4131
rect 38936 4088 38988 4097
rect 43536 4131 43588 4140
rect 43536 4097 43545 4131
rect 43545 4097 43579 4131
rect 43579 4097 43588 4131
rect 43536 4088 43588 4097
rect 46112 4156 46164 4208
rect 55404 4156 55456 4208
rect 55496 4156 55548 4208
rect 68100 4156 68152 4208
rect 47952 4088 48004 4140
rect 53288 4088 53340 4140
rect 55864 4088 55916 4140
rect 37188 3952 37240 4004
rect 42248 4020 42300 4072
rect 43352 4020 43404 4072
rect 45468 4063 45520 4072
rect 45468 4029 45477 4063
rect 45477 4029 45511 4063
rect 45511 4029 45520 4063
rect 45468 4020 45520 4029
rect 41328 3952 41380 4004
rect 47584 4020 47636 4072
rect 47768 4020 47820 4072
rect 49332 4020 49384 4072
rect 49424 4020 49476 4072
rect 51540 3952 51592 4004
rect 52276 3952 52328 4004
rect 58624 3952 58676 4004
rect 25228 3927 25280 3936
rect 25228 3893 25237 3927
rect 25237 3893 25271 3927
rect 25271 3893 25280 3927
rect 25228 3884 25280 3893
rect 25320 3927 25372 3936
rect 25320 3893 25329 3927
rect 25329 3893 25363 3927
rect 25363 3893 25372 3927
rect 25320 3884 25372 3893
rect 26056 3927 26108 3936
rect 26056 3893 26065 3927
rect 26065 3893 26099 3927
rect 26099 3893 26108 3927
rect 26056 3884 26108 3893
rect 28448 3884 28500 3936
rect 29000 3884 29052 3936
rect 29092 3884 29144 3936
rect 30932 3884 30984 3936
rect 31208 3927 31260 3936
rect 31208 3893 31217 3927
rect 31217 3893 31251 3927
rect 31251 3893 31260 3927
rect 31208 3884 31260 3893
rect 32864 3927 32916 3936
rect 32864 3893 32873 3927
rect 32873 3893 32907 3927
rect 32907 3893 32916 3927
rect 32864 3884 32916 3893
rect 33232 3884 33284 3936
rect 34060 3884 34112 3936
rect 35072 3927 35124 3936
rect 35072 3893 35081 3927
rect 35081 3893 35115 3927
rect 35115 3893 35124 3927
rect 35072 3884 35124 3893
rect 36820 3884 36872 3936
rect 41512 3927 41564 3936
rect 41512 3893 41521 3927
rect 41521 3893 41555 3927
rect 41555 3893 41564 3927
rect 41512 3884 41564 3893
rect 43812 3884 43864 3936
rect 50804 3884 50856 3936
rect 55864 3884 55916 3936
rect 65248 3884 65300 3936
rect 1858 3782 1910 3834
rect 1922 3782 1974 3834
rect 1986 3782 2038 3834
rect 2050 3782 2102 3834
rect 2114 3782 2166 3834
rect 11858 3782 11910 3834
rect 11922 3782 11974 3834
rect 11986 3782 12038 3834
rect 12050 3782 12102 3834
rect 12114 3782 12166 3834
rect 21858 3782 21910 3834
rect 21922 3782 21974 3834
rect 21986 3782 22038 3834
rect 22050 3782 22102 3834
rect 22114 3782 22166 3834
rect 31858 3782 31910 3834
rect 31922 3782 31974 3834
rect 31986 3782 32038 3834
rect 32050 3782 32102 3834
rect 32114 3782 32166 3834
rect 41858 3782 41910 3834
rect 41922 3782 41974 3834
rect 41986 3782 42038 3834
rect 42050 3782 42102 3834
rect 42114 3782 42166 3834
rect 51858 3782 51910 3834
rect 51922 3782 51974 3834
rect 51986 3782 52038 3834
rect 52050 3782 52102 3834
rect 52114 3782 52166 3834
rect 61858 3782 61910 3834
rect 61922 3782 61974 3834
rect 61986 3782 62038 3834
rect 62050 3782 62102 3834
rect 62114 3782 62166 3834
rect 71858 3782 71910 3834
rect 71922 3782 71974 3834
rect 71986 3782 72038 3834
rect 72050 3782 72102 3834
rect 72114 3782 72166 3834
rect 23664 3476 23716 3528
rect 25320 3476 25372 3528
rect 27896 3680 27948 3732
rect 29828 3680 29880 3732
rect 29920 3680 29972 3732
rect 30748 3680 30800 3732
rect 33416 3680 33468 3732
rect 35256 3680 35308 3732
rect 27344 3544 27396 3596
rect 26424 3519 26476 3528
rect 26424 3485 26433 3519
rect 26433 3485 26467 3519
rect 26467 3485 26476 3519
rect 26424 3476 26476 3485
rect 29736 3612 29788 3664
rect 40132 3680 40184 3732
rect 27896 3544 27948 3596
rect 29092 3544 29144 3596
rect 27804 3519 27856 3528
rect 27804 3485 27813 3519
rect 27813 3485 27847 3519
rect 27847 3485 27856 3519
rect 27804 3476 27856 3485
rect 27988 3519 28040 3528
rect 27988 3485 27997 3519
rect 27997 3485 28031 3519
rect 28031 3485 28040 3519
rect 27988 3476 28040 3485
rect 32864 3544 32916 3596
rect 34060 3544 34112 3596
rect 40868 3655 40920 3664
rect 40868 3621 40877 3655
rect 40877 3621 40911 3655
rect 40911 3621 40920 3655
rect 40868 3612 40920 3621
rect 42248 3680 42300 3732
rect 43352 3680 43404 3732
rect 45008 3612 45060 3664
rect 41512 3544 41564 3596
rect 42248 3544 42300 3596
rect 44732 3544 44784 3596
rect 26608 3408 26660 3460
rect 30564 3408 30616 3460
rect 24032 3340 24084 3392
rect 24952 3383 25004 3392
rect 24952 3349 24961 3383
rect 24961 3349 24995 3383
rect 24995 3349 25004 3383
rect 24952 3340 25004 3349
rect 26976 3340 27028 3392
rect 27068 3383 27120 3392
rect 27068 3349 27077 3383
rect 27077 3349 27111 3383
rect 27111 3349 27120 3383
rect 27068 3340 27120 3349
rect 29184 3340 29236 3392
rect 30104 3383 30156 3392
rect 30104 3349 30113 3383
rect 30113 3349 30147 3383
rect 30147 3349 30156 3383
rect 30104 3340 30156 3349
rect 30748 3408 30800 3460
rect 31668 3340 31720 3392
rect 32312 3519 32364 3528
rect 32312 3485 32321 3519
rect 32321 3485 32355 3519
rect 32355 3485 32364 3519
rect 32312 3476 32364 3485
rect 32588 3476 32640 3528
rect 34704 3519 34756 3528
rect 34704 3485 34713 3519
rect 34713 3485 34747 3519
rect 34747 3485 34756 3519
rect 34704 3476 34756 3485
rect 35900 3476 35952 3528
rect 36084 3476 36136 3528
rect 38384 3519 38436 3528
rect 38384 3485 38393 3519
rect 38393 3485 38427 3519
rect 38427 3485 38436 3519
rect 38384 3476 38436 3485
rect 39120 3519 39172 3528
rect 39120 3485 39129 3519
rect 39129 3485 39163 3519
rect 39163 3485 39172 3519
rect 39120 3476 39172 3485
rect 40316 3519 40368 3528
rect 40316 3485 40325 3519
rect 40325 3485 40359 3519
rect 40359 3485 40368 3519
rect 40316 3476 40368 3485
rect 40592 3519 40644 3528
rect 40592 3485 40601 3519
rect 40601 3485 40635 3519
rect 40635 3485 40644 3519
rect 40592 3476 40644 3485
rect 41328 3519 41380 3528
rect 41328 3485 41337 3519
rect 41337 3485 41371 3519
rect 41371 3485 41380 3519
rect 41328 3476 41380 3485
rect 41604 3476 41656 3528
rect 44640 3519 44692 3528
rect 44640 3485 44649 3519
rect 44649 3485 44683 3519
rect 44683 3485 44692 3519
rect 44640 3476 44692 3485
rect 45560 3476 45612 3528
rect 48412 3680 48464 3732
rect 49424 3723 49476 3732
rect 49424 3689 49433 3723
rect 49433 3689 49467 3723
rect 49467 3689 49476 3723
rect 49424 3680 49476 3689
rect 49608 3680 49660 3732
rect 55864 3680 55916 3732
rect 48320 3612 48372 3664
rect 54668 3612 54720 3664
rect 65524 3680 65576 3732
rect 59084 3612 59136 3664
rect 63592 3612 63644 3664
rect 49884 3544 49936 3596
rect 53932 3544 53984 3596
rect 64696 3612 64748 3664
rect 33140 3408 33192 3460
rect 32772 3340 32824 3392
rect 32956 3383 33008 3392
rect 32956 3349 32965 3383
rect 32965 3349 32999 3383
rect 32999 3349 33008 3383
rect 32956 3340 33008 3349
rect 33048 3340 33100 3392
rect 35164 3408 35216 3460
rect 35624 3408 35676 3460
rect 42340 3408 42392 3460
rect 47492 3476 47544 3528
rect 48964 3476 49016 3528
rect 47124 3408 47176 3460
rect 50712 3519 50764 3528
rect 50712 3485 50721 3519
rect 50721 3485 50755 3519
rect 50755 3485 50764 3519
rect 50712 3476 50764 3485
rect 52644 3476 52696 3528
rect 53012 3519 53064 3528
rect 53012 3485 53021 3519
rect 53021 3485 53055 3519
rect 53055 3485 53064 3519
rect 53012 3476 53064 3485
rect 55956 3476 56008 3528
rect 60372 3476 60424 3528
rect 51540 3408 51592 3460
rect 54024 3408 54076 3460
rect 59176 3408 59228 3460
rect 33692 3383 33744 3392
rect 33692 3349 33701 3383
rect 33701 3349 33735 3383
rect 33735 3349 33744 3383
rect 33692 3340 33744 3349
rect 33784 3383 33836 3392
rect 33784 3349 33793 3383
rect 33793 3349 33827 3383
rect 33827 3349 33836 3383
rect 33784 3340 33836 3349
rect 34888 3340 34940 3392
rect 37464 3340 37516 3392
rect 42524 3340 42576 3392
rect 43444 3340 43496 3392
rect 43536 3340 43588 3392
rect 45468 3340 45520 3392
rect 46940 3340 46992 3392
rect 47032 3383 47084 3392
rect 47032 3349 47041 3383
rect 47041 3349 47075 3383
rect 47075 3349 47084 3383
rect 47032 3340 47084 3349
rect 49976 3340 50028 3392
rect 50436 3340 50488 3392
rect 51448 3383 51500 3392
rect 51448 3349 51457 3383
rect 51457 3349 51491 3383
rect 51491 3349 51500 3383
rect 51448 3340 51500 3349
rect 52368 3383 52420 3392
rect 52368 3349 52377 3383
rect 52377 3349 52411 3383
rect 52411 3349 52420 3383
rect 52368 3340 52420 3349
rect 55588 3340 55640 3392
rect 58164 3383 58216 3392
rect 58164 3349 58173 3383
rect 58173 3349 58207 3383
rect 58207 3349 58216 3383
rect 58164 3340 58216 3349
rect 60740 3408 60792 3460
rect 64696 3476 64748 3528
rect 64972 3476 65024 3528
rect 72424 3476 72476 3528
rect 70584 3408 70636 3460
rect 72516 3340 72568 3392
rect 4210 3238 4262 3290
rect 4274 3238 4326 3290
rect 4338 3238 4390 3290
rect 4402 3238 4454 3290
rect 4466 3238 4518 3290
rect 14210 3238 14262 3290
rect 14274 3238 14326 3290
rect 14338 3238 14390 3290
rect 14402 3238 14454 3290
rect 14466 3238 14518 3290
rect 24210 3238 24262 3290
rect 24274 3238 24326 3290
rect 24338 3238 24390 3290
rect 24402 3238 24454 3290
rect 24466 3238 24518 3290
rect 34210 3238 34262 3290
rect 34274 3238 34326 3290
rect 34338 3238 34390 3290
rect 34402 3238 34454 3290
rect 34466 3238 34518 3290
rect 44210 3238 44262 3290
rect 44274 3238 44326 3290
rect 44338 3238 44390 3290
rect 44402 3238 44454 3290
rect 44466 3238 44518 3290
rect 54210 3238 54262 3290
rect 54274 3238 54326 3290
rect 54338 3238 54390 3290
rect 54402 3238 54454 3290
rect 54466 3238 54518 3290
rect 64210 3238 64262 3290
rect 64274 3238 64326 3290
rect 64338 3238 64390 3290
rect 64402 3238 64454 3290
rect 64466 3238 64518 3290
rect 74210 3238 74262 3290
rect 74274 3238 74326 3290
rect 74338 3238 74390 3290
rect 74402 3238 74454 3290
rect 74466 3238 74518 3290
rect 24584 3136 24636 3188
rect 27068 3136 27120 3188
rect 25964 3068 26016 3120
rect 27620 3068 27672 3120
rect 29184 3068 29236 3120
rect 25044 3000 25096 3052
rect 32220 3136 32272 3188
rect 32496 3136 32548 3188
rect 32588 3179 32640 3188
rect 32588 3145 32597 3179
rect 32597 3145 32631 3179
rect 32631 3145 32640 3179
rect 32588 3136 32640 3145
rect 34980 3136 35032 3188
rect 35992 3136 36044 3188
rect 36360 3136 36412 3188
rect 38016 3179 38068 3188
rect 38016 3145 38025 3179
rect 38025 3145 38059 3179
rect 38059 3145 38068 3179
rect 38016 3136 38068 3145
rect 22376 2975 22428 2984
rect 22376 2941 22385 2975
rect 22385 2941 22419 2975
rect 22419 2941 22428 2975
rect 22376 2932 22428 2941
rect 23112 2975 23164 2984
rect 23112 2941 23121 2975
rect 23121 2941 23155 2975
rect 23155 2941 23164 2975
rect 23112 2932 23164 2941
rect 23848 2975 23900 2984
rect 23848 2941 23857 2975
rect 23857 2941 23891 2975
rect 23891 2941 23900 2975
rect 23848 2932 23900 2941
rect 25320 2975 25372 2984
rect 25320 2941 25329 2975
rect 25329 2941 25363 2975
rect 25363 2941 25372 2975
rect 25320 2932 25372 2941
rect 20996 2864 21048 2916
rect 23572 2864 23624 2916
rect 27160 2975 27212 2984
rect 27160 2941 27169 2975
rect 27169 2941 27203 2975
rect 27203 2941 27212 2975
rect 27160 2932 27212 2941
rect 27896 2932 27948 2984
rect 29828 3000 29880 3052
rect 29276 2932 29328 2984
rect 22284 2796 22336 2848
rect 23480 2796 23532 2848
rect 24584 2839 24636 2848
rect 24584 2805 24593 2839
rect 24593 2805 24627 2839
rect 24627 2805 24636 2839
rect 24584 2796 24636 2805
rect 25412 2796 25464 2848
rect 28172 2864 28224 2916
rect 30472 2975 30524 2984
rect 30472 2941 30481 2975
rect 30481 2941 30515 2975
rect 30515 2941 30524 2975
rect 30472 2932 30524 2941
rect 31208 3043 31260 3052
rect 31208 3009 31217 3043
rect 31217 3009 31251 3043
rect 31251 3009 31260 3043
rect 31208 3000 31260 3009
rect 33048 3000 33100 3052
rect 33232 3043 33284 3052
rect 33232 3009 33241 3043
rect 33241 3009 33275 3043
rect 33275 3009 33284 3043
rect 33232 3000 33284 3009
rect 33692 3000 33744 3052
rect 40224 3068 40276 3120
rect 42340 3179 42392 3188
rect 42340 3145 42349 3179
rect 42349 3145 42383 3179
rect 42383 3145 42392 3179
rect 42340 3136 42392 3145
rect 44640 3136 44692 3188
rect 43536 3068 43588 3120
rect 47492 3179 47544 3188
rect 47492 3145 47501 3179
rect 47501 3145 47535 3179
rect 47535 3145 47544 3179
rect 47492 3136 47544 3145
rect 48964 3179 49016 3188
rect 48964 3145 48973 3179
rect 48973 3145 49007 3179
rect 49007 3145 49016 3179
rect 48964 3136 49016 3145
rect 51356 3068 51408 3120
rect 52368 3068 52420 3120
rect 52644 3179 52696 3188
rect 52644 3145 52653 3179
rect 52653 3145 52687 3179
rect 52687 3145 52696 3179
rect 52644 3136 52696 3145
rect 53840 3068 53892 3120
rect 59268 3068 59320 3120
rect 34888 3043 34940 3052
rect 34888 3009 34897 3043
rect 34897 3009 34931 3043
rect 34931 3009 34940 3043
rect 34888 3000 34940 3009
rect 35624 3043 35676 3052
rect 35624 3009 35633 3043
rect 35633 3009 35667 3043
rect 35667 3009 35676 3043
rect 35624 3000 35676 3009
rect 36820 3043 36872 3052
rect 36820 3009 36829 3043
rect 36829 3009 36863 3043
rect 36863 3009 36872 3043
rect 36820 3000 36872 3009
rect 39856 3043 39908 3052
rect 39856 3009 39865 3043
rect 39865 3009 39899 3043
rect 39899 3009 39908 3043
rect 39856 3000 39908 3009
rect 40040 3000 40092 3052
rect 34980 2932 35032 2984
rect 37280 2975 37332 2984
rect 37280 2941 37289 2975
rect 37289 2941 37323 2975
rect 37323 2941 37332 2975
rect 37280 2932 37332 2941
rect 40132 2932 40184 2984
rect 40224 2975 40276 2984
rect 40224 2941 40233 2975
rect 40233 2941 40267 2975
rect 40267 2941 40276 2975
rect 40224 2932 40276 2941
rect 41696 2864 41748 2916
rect 43812 3043 43864 3052
rect 43812 3009 43821 3043
rect 43821 3009 43855 3043
rect 43855 3009 43864 3043
rect 43812 3000 43864 3009
rect 48872 3000 48924 3052
rect 50436 3043 50488 3052
rect 50436 3009 50445 3043
rect 50445 3009 50479 3043
rect 50479 3009 50488 3043
rect 50436 3000 50488 3009
rect 51724 3000 51776 3052
rect 54944 3000 54996 3052
rect 55588 3043 55640 3052
rect 55588 3009 55597 3043
rect 55597 3009 55631 3043
rect 55631 3009 55640 3043
rect 55588 3000 55640 3009
rect 58164 3000 58216 3052
rect 59176 3043 59228 3052
rect 59176 3009 59185 3043
rect 59185 3009 59219 3043
rect 59219 3009 59228 3043
rect 59176 3000 59228 3009
rect 60740 3179 60792 3188
rect 60740 3145 60749 3179
rect 60749 3145 60783 3179
rect 60783 3145 60792 3179
rect 60740 3136 60792 3145
rect 70952 3136 71004 3188
rect 64972 3068 65024 3120
rect 68376 3068 68428 3120
rect 63408 3000 63460 3052
rect 66812 3000 66864 3052
rect 69112 3000 69164 3052
rect 72700 3000 72752 3052
rect 42984 2975 43036 2984
rect 42984 2941 42993 2975
rect 42993 2941 43027 2975
rect 43027 2941 43036 2975
rect 42984 2932 43036 2941
rect 44640 2975 44692 2984
rect 44640 2941 44649 2975
rect 44649 2941 44683 2975
rect 44683 2941 44692 2975
rect 44640 2932 44692 2941
rect 46112 2975 46164 2984
rect 46112 2941 46121 2975
rect 46121 2941 46155 2975
rect 46155 2941 46164 2975
rect 46112 2932 46164 2941
rect 46848 2932 46900 2984
rect 45376 2864 45428 2916
rect 46020 2864 46072 2916
rect 48780 2975 48832 2984
rect 48780 2941 48789 2975
rect 48789 2941 48823 2975
rect 48823 2941 48832 2975
rect 48780 2932 48832 2941
rect 49332 2932 49384 2984
rect 27528 2796 27580 2848
rect 28080 2796 28132 2848
rect 30012 2796 30064 2848
rect 33968 2796 34020 2848
rect 36176 2839 36228 2848
rect 36176 2805 36185 2839
rect 36185 2805 36219 2839
rect 36219 2805 36228 2839
rect 36176 2796 36228 2805
rect 38752 2839 38804 2848
rect 38752 2805 38761 2839
rect 38761 2805 38795 2839
rect 38795 2805 38804 2839
rect 38752 2796 38804 2805
rect 41420 2796 41472 2848
rect 41512 2839 41564 2848
rect 41512 2805 41521 2839
rect 41521 2805 41555 2839
rect 41555 2805 41564 2839
rect 41512 2796 41564 2805
rect 42340 2796 42392 2848
rect 45928 2796 45980 2848
rect 47400 2796 47452 2848
rect 51632 2932 51684 2984
rect 52644 2932 52696 2984
rect 54576 2932 54628 2984
rect 55680 2932 55732 2984
rect 57060 2932 57112 2984
rect 59820 2932 59872 2984
rect 61384 2975 61436 2984
rect 61384 2941 61393 2975
rect 61393 2941 61427 2975
rect 61427 2941 61436 2975
rect 61384 2932 61436 2941
rect 61568 2975 61620 2984
rect 61568 2941 61577 2975
rect 61577 2941 61611 2975
rect 61611 2941 61620 2975
rect 61568 2932 61620 2941
rect 63316 2932 63368 2984
rect 65248 2975 65300 2984
rect 65248 2941 65257 2975
rect 65257 2941 65291 2975
rect 65291 2941 65300 2975
rect 65248 2932 65300 2941
rect 51356 2864 51408 2916
rect 52920 2864 52972 2916
rect 55312 2864 55364 2916
rect 56600 2864 56652 2916
rect 58532 2864 58584 2916
rect 62580 2864 62632 2916
rect 51080 2839 51132 2848
rect 51080 2805 51089 2839
rect 51089 2805 51123 2839
rect 51123 2805 51132 2839
rect 51080 2796 51132 2805
rect 51172 2839 51224 2848
rect 51172 2805 51181 2839
rect 51181 2805 51215 2839
rect 51215 2805 51224 2839
rect 51172 2796 51224 2805
rect 55220 2796 55272 2848
rect 56876 2796 56928 2848
rect 56968 2839 57020 2848
rect 56968 2805 56977 2839
rect 56977 2805 57011 2839
rect 57011 2805 57020 2839
rect 56968 2796 57020 2805
rect 58900 2796 58952 2848
rect 59912 2839 59964 2848
rect 59912 2805 59921 2839
rect 59921 2805 59955 2839
rect 59955 2805 59964 2839
rect 59912 2796 59964 2805
rect 61108 2796 61160 2848
rect 64972 2796 65024 2848
rect 69020 2975 69072 2984
rect 69020 2941 69029 2975
rect 69029 2941 69063 2975
rect 69063 2941 69072 2975
rect 69020 2932 69072 2941
rect 69480 2932 69532 2984
rect 71044 2975 71096 2984
rect 71044 2941 71053 2975
rect 71053 2941 71087 2975
rect 71087 2941 71096 2975
rect 71044 2932 71096 2941
rect 73252 2932 73304 2984
rect 69388 2864 69440 2916
rect 70676 2864 70728 2916
rect 66260 2796 66312 2848
rect 66996 2839 67048 2848
rect 66996 2805 67005 2839
rect 67005 2805 67039 2839
rect 67039 2805 67048 2839
rect 66996 2796 67048 2805
rect 68468 2796 68520 2848
rect 70860 2796 70912 2848
rect 72240 2796 72292 2848
rect 1858 2694 1910 2746
rect 1922 2694 1974 2746
rect 1986 2694 2038 2746
rect 2050 2694 2102 2746
rect 2114 2694 2166 2746
rect 11858 2694 11910 2746
rect 11922 2694 11974 2746
rect 11986 2694 12038 2746
rect 12050 2694 12102 2746
rect 12114 2694 12166 2746
rect 21858 2694 21910 2746
rect 21922 2694 21974 2746
rect 21986 2694 22038 2746
rect 22050 2694 22102 2746
rect 22114 2694 22166 2746
rect 31858 2694 31910 2746
rect 31922 2694 31974 2746
rect 31986 2694 32038 2746
rect 32050 2694 32102 2746
rect 32114 2694 32166 2746
rect 41858 2694 41910 2746
rect 41922 2694 41974 2746
rect 41986 2694 42038 2746
rect 42050 2694 42102 2746
rect 42114 2694 42166 2746
rect 51858 2694 51910 2746
rect 51922 2694 51974 2746
rect 51986 2694 52038 2746
rect 52050 2694 52102 2746
rect 52114 2694 52166 2746
rect 61858 2694 61910 2746
rect 61922 2694 61974 2746
rect 61986 2694 62038 2746
rect 62050 2694 62102 2746
rect 62114 2694 62166 2746
rect 71858 2694 71910 2746
rect 71922 2694 71974 2746
rect 71986 2694 72038 2746
rect 72050 2694 72102 2746
rect 72114 2694 72166 2746
rect 23112 2592 23164 2644
rect 23848 2592 23900 2644
rect 24032 2524 24084 2576
rect 24032 2388 24084 2440
rect 27712 2592 27764 2644
rect 27988 2592 28040 2644
rect 29368 2592 29420 2644
rect 29552 2592 29604 2644
rect 30472 2592 30524 2644
rect 32312 2592 32364 2644
rect 34612 2592 34664 2644
rect 36084 2592 36136 2644
rect 36912 2635 36964 2644
rect 36912 2601 36921 2635
rect 36921 2601 36955 2635
rect 36955 2601 36964 2635
rect 36912 2592 36964 2601
rect 38384 2592 38436 2644
rect 40224 2592 40276 2644
rect 42984 2592 43036 2644
rect 44640 2592 44692 2644
rect 45560 2592 45612 2644
rect 46112 2592 46164 2644
rect 48780 2592 48832 2644
rect 49516 2592 49568 2644
rect 50712 2592 50764 2644
rect 51540 2635 51592 2644
rect 51540 2601 51549 2635
rect 51549 2601 51583 2635
rect 51583 2601 51592 2635
rect 51540 2592 51592 2601
rect 53012 2635 53064 2644
rect 53012 2601 53021 2635
rect 53021 2601 53055 2635
rect 53055 2601 53064 2635
rect 53012 2592 53064 2601
rect 26608 2524 26660 2576
rect 30012 2567 30064 2576
rect 30012 2533 30021 2567
rect 30021 2533 30055 2567
rect 30055 2533 30064 2567
rect 30012 2524 30064 2533
rect 32680 2524 32732 2576
rect 34704 2524 34756 2576
rect 34796 2524 34848 2576
rect 54668 2524 54720 2576
rect 55956 2567 56008 2576
rect 55956 2533 55965 2567
rect 55965 2533 55999 2567
rect 55999 2533 56008 2567
rect 55956 2524 56008 2533
rect 60648 2524 60700 2576
rect 61568 2524 61620 2576
rect 63316 2567 63368 2576
rect 63316 2533 63325 2567
rect 63325 2533 63359 2567
rect 63359 2533 63368 2567
rect 63316 2524 63368 2533
rect 64696 2524 64748 2576
rect 65248 2592 65300 2644
rect 66260 2635 66312 2644
rect 66260 2601 66269 2635
rect 66269 2601 66303 2635
rect 66303 2601 66312 2635
rect 66260 2592 66312 2601
rect 69112 2635 69164 2644
rect 69112 2601 69121 2635
rect 69121 2601 69155 2635
rect 69155 2601 69164 2635
rect 69112 2592 69164 2601
rect 71044 2592 71096 2644
rect 69664 2524 69716 2576
rect 30104 2456 30156 2508
rect 30748 2499 30800 2508
rect 30748 2465 30757 2499
rect 30757 2465 30791 2499
rect 30791 2465 30800 2499
rect 30748 2456 30800 2465
rect 31116 2456 31168 2508
rect 32404 2456 32456 2508
rect 33784 2499 33836 2508
rect 33784 2465 33793 2499
rect 33793 2465 33827 2499
rect 33827 2465 33836 2499
rect 33784 2456 33836 2465
rect 24584 2320 24636 2372
rect 25412 2431 25464 2440
rect 25412 2397 25421 2431
rect 25421 2397 25455 2431
rect 25455 2397 25464 2431
rect 25412 2388 25464 2397
rect 27068 2388 27120 2440
rect 28264 2388 28316 2440
rect 28448 2431 28500 2440
rect 28448 2397 28457 2431
rect 28457 2397 28491 2431
rect 28491 2397 28500 2431
rect 28448 2388 28500 2397
rect 31024 2388 31076 2440
rect 26792 2320 26844 2372
rect 27528 2320 27580 2372
rect 28908 2320 28960 2372
rect 33048 2431 33100 2440
rect 33048 2397 33057 2431
rect 33057 2397 33091 2431
rect 33091 2397 33100 2431
rect 33048 2388 33100 2397
rect 35532 2431 35584 2440
rect 35532 2397 35541 2431
rect 35541 2397 35575 2431
rect 35575 2397 35584 2431
rect 35532 2388 35584 2397
rect 36176 2456 36228 2508
rect 37832 2456 37884 2508
rect 38752 2499 38804 2508
rect 38752 2465 38761 2499
rect 38761 2465 38795 2499
rect 38795 2465 38804 2499
rect 38752 2456 38804 2465
rect 41512 2456 41564 2508
rect 42524 2456 42576 2508
rect 43444 2499 43496 2508
rect 43444 2465 43453 2499
rect 43453 2465 43487 2499
rect 43487 2465 43496 2499
rect 43444 2456 43496 2465
rect 46940 2499 46992 2508
rect 46940 2465 46949 2499
rect 46949 2465 46983 2499
rect 46983 2465 46992 2499
rect 46940 2456 46992 2465
rect 47124 2499 47176 2508
rect 47124 2465 47133 2499
rect 47133 2465 47167 2499
rect 47167 2465 47176 2499
rect 47124 2456 47176 2465
rect 47308 2456 47360 2508
rect 49792 2456 49844 2508
rect 49976 2456 50028 2508
rect 51080 2456 51132 2508
rect 54024 2456 54076 2508
rect 55220 2499 55272 2508
rect 55220 2465 55229 2499
rect 55229 2465 55263 2499
rect 55263 2465 55272 2499
rect 55220 2456 55272 2465
rect 56600 2499 56652 2508
rect 56600 2465 56609 2499
rect 56609 2465 56643 2499
rect 56643 2465 56652 2499
rect 56600 2456 56652 2465
rect 56876 2456 56928 2508
rect 58900 2499 58952 2508
rect 58900 2465 58909 2499
rect 58909 2465 58943 2499
rect 58943 2465 58952 2499
rect 58900 2456 58952 2465
rect 59912 2456 59964 2508
rect 61108 2499 61160 2508
rect 61108 2465 61117 2499
rect 61117 2465 61151 2499
rect 61151 2465 61160 2499
rect 61108 2456 61160 2465
rect 36360 2388 36412 2440
rect 37648 2388 37700 2440
rect 34612 2320 34664 2372
rect 36268 2320 36320 2372
rect 41052 2431 41104 2440
rect 41052 2397 41061 2431
rect 41061 2397 41095 2431
rect 41095 2397 41104 2431
rect 41052 2388 41104 2397
rect 40776 2320 40828 2372
rect 45560 2431 45612 2440
rect 45560 2397 45569 2431
rect 45569 2397 45603 2431
rect 45603 2397 45612 2431
rect 45560 2388 45612 2397
rect 46112 2388 46164 2440
rect 49424 2388 49476 2440
rect 51356 2431 51408 2440
rect 51356 2397 51365 2431
rect 51365 2397 51399 2431
rect 51399 2397 51408 2431
rect 51356 2388 51408 2397
rect 51448 2388 51500 2440
rect 56692 2388 56744 2440
rect 58440 2388 58492 2440
rect 59728 2388 59780 2440
rect 61568 2388 61620 2440
rect 47216 2320 47268 2372
rect 47676 2320 47728 2372
rect 50160 2320 50212 2372
rect 57244 2320 57296 2372
rect 61660 2320 61712 2372
rect 62580 2499 62632 2508
rect 62580 2465 62589 2499
rect 62589 2465 62623 2499
rect 62623 2465 62632 2499
rect 62580 2456 62632 2465
rect 62672 2456 62724 2508
rect 62764 2388 62816 2440
rect 64788 2320 64840 2372
rect 64972 2499 65024 2508
rect 64972 2465 64981 2499
rect 64981 2465 65015 2499
rect 65015 2465 65024 2499
rect 64972 2456 65024 2465
rect 66996 2499 67048 2508
rect 66996 2465 67005 2499
rect 67005 2465 67039 2499
rect 67039 2465 67048 2499
rect 66996 2456 67048 2465
rect 68468 2499 68520 2508
rect 68468 2465 68477 2499
rect 68477 2465 68511 2499
rect 68511 2465 68520 2499
rect 68468 2456 68520 2465
rect 65340 2388 65392 2440
rect 66076 2431 66128 2440
rect 66076 2397 66085 2431
rect 66085 2397 66119 2431
rect 66119 2397 66128 2431
rect 66076 2388 66128 2397
rect 67088 2388 67140 2440
rect 68376 2388 68428 2440
rect 71228 2524 71280 2576
rect 70124 2499 70176 2508
rect 70124 2465 70133 2499
rect 70133 2465 70167 2499
rect 70167 2465 70176 2499
rect 70124 2456 70176 2465
rect 70676 2499 70728 2508
rect 70676 2465 70685 2499
rect 70685 2465 70719 2499
rect 70719 2465 70728 2499
rect 70676 2456 70728 2465
rect 72240 2499 72292 2508
rect 72240 2465 72249 2499
rect 72249 2465 72283 2499
rect 72283 2465 72292 2499
rect 72240 2456 72292 2465
rect 72240 2320 72292 2372
rect 23480 2295 23532 2304
rect 23480 2261 23489 2295
rect 23489 2261 23523 2295
rect 23523 2261 23532 2295
rect 23480 2252 23532 2261
rect 25320 2252 25372 2304
rect 28632 2252 28684 2304
rect 34888 2252 34940 2304
rect 35716 2252 35768 2304
rect 39580 2252 39632 2304
rect 40316 2252 40368 2304
rect 44824 2252 44876 2304
rect 44916 2252 44968 2304
rect 46940 2252 46992 2304
rect 48504 2295 48556 2304
rect 48504 2261 48513 2295
rect 48513 2261 48547 2295
rect 48547 2261 48556 2295
rect 48504 2252 48556 2261
rect 53196 2252 53248 2304
rect 56048 2252 56100 2304
rect 59452 2252 59504 2304
rect 59544 2295 59596 2304
rect 59544 2261 59553 2295
rect 59553 2261 59587 2295
rect 59587 2261 59596 2295
rect 59544 2252 59596 2261
rect 61200 2252 61252 2304
rect 62488 2252 62540 2304
rect 64972 2252 65024 2304
rect 68100 2252 68152 2304
rect 69756 2252 69808 2304
rect 70676 2252 70728 2304
rect 74632 2252 74684 2304
rect 4210 2150 4262 2202
rect 4274 2150 4326 2202
rect 4338 2150 4390 2202
rect 4402 2150 4454 2202
rect 4466 2150 4518 2202
rect 14210 2150 14262 2202
rect 14274 2150 14326 2202
rect 14338 2150 14390 2202
rect 14402 2150 14454 2202
rect 14466 2150 14518 2202
rect 24210 2150 24262 2202
rect 24274 2150 24326 2202
rect 24338 2150 24390 2202
rect 24402 2150 24454 2202
rect 24466 2150 24518 2202
rect 34210 2150 34262 2202
rect 34274 2150 34326 2202
rect 34338 2150 34390 2202
rect 34402 2150 34454 2202
rect 34466 2150 34518 2202
rect 44210 2150 44262 2202
rect 44274 2150 44326 2202
rect 44338 2150 44390 2202
rect 44402 2150 44454 2202
rect 44466 2150 44518 2202
rect 54210 2150 54262 2202
rect 54274 2150 54326 2202
rect 54338 2150 54390 2202
rect 54402 2150 54454 2202
rect 54466 2150 54518 2202
rect 64210 2150 64262 2202
rect 64274 2150 64326 2202
rect 64338 2150 64390 2202
rect 64402 2150 64454 2202
rect 64466 2150 64518 2202
rect 74210 2150 74262 2202
rect 74274 2150 74326 2202
rect 74338 2150 74390 2202
rect 74402 2150 74454 2202
rect 74466 2150 74518 2202
rect 22376 2048 22428 2100
rect 24952 2048 25004 2100
rect 26240 2048 26292 2100
rect 27620 2048 27672 2100
rect 23480 1955 23532 1964
rect 23480 1921 23489 1955
rect 23489 1921 23523 1955
rect 23523 1921 23532 1955
rect 23480 1912 23532 1921
rect 25228 1912 25280 1964
rect 26884 1955 26936 1964
rect 26884 1921 26893 1955
rect 26893 1921 26927 1955
rect 26927 1921 26936 1955
rect 26884 1912 26936 1921
rect 26976 1912 27028 1964
rect 29000 1955 29052 1964
rect 29000 1921 29009 1955
rect 29009 1921 29043 1955
rect 29043 1921 29052 1955
rect 29000 1912 29052 1921
rect 33324 2048 33376 2100
rect 36268 2091 36320 2100
rect 36268 2057 36277 2091
rect 36277 2057 36311 2091
rect 36311 2057 36320 2091
rect 36268 2048 36320 2057
rect 37280 2048 37332 2100
rect 39120 2048 39172 2100
rect 39856 2048 39908 2100
rect 40592 2048 40644 2100
rect 45376 2091 45428 2100
rect 45376 2057 45385 2091
rect 45385 2057 45419 2091
rect 45419 2057 45428 2091
rect 45376 2048 45428 2057
rect 46112 2091 46164 2100
rect 46112 2057 46121 2091
rect 46121 2057 46155 2091
rect 46155 2057 46164 2091
rect 46112 2048 46164 2057
rect 23572 1887 23624 1896
rect 23572 1853 23581 1887
rect 23581 1853 23615 1887
rect 23615 1853 23624 1887
rect 23572 1844 23624 1853
rect 24032 1844 24084 1896
rect 25320 1844 25372 1896
rect 25596 1844 25648 1896
rect 26148 1887 26200 1896
rect 26148 1853 26157 1887
rect 26157 1853 26191 1887
rect 26191 1853 26200 1887
rect 26148 1844 26200 1853
rect 36544 1980 36596 2032
rect 55864 2048 55916 2100
rect 56508 2048 56560 2100
rect 58440 2091 58492 2100
rect 58440 2057 58449 2091
rect 58449 2057 58483 2091
rect 58483 2057 58492 2091
rect 58440 2048 58492 2057
rect 60372 2048 60424 2100
rect 61384 2048 61436 2100
rect 66076 2091 66128 2100
rect 66076 2057 66085 2091
rect 66085 2057 66119 2091
rect 66119 2057 66128 2091
rect 66076 2048 66128 2057
rect 69020 2048 69072 2100
rect 32864 1912 32916 1964
rect 34796 1912 34848 1964
rect 35624 1912 35676 1964
rect 35716 1955 35768 1964
rect 35716 1921 35725 1955
rect 35725 1921 35759 1955
rect 35759 1921 35768 1955
rect 35716 1912 35768 1921
rect 37464 1912 37516 1964
rect 39580 1955 39632 1964
rect 39580 1921 39589 1955
rect 39589 1921 39623 1955
rect 39623 1921 39632 1955
rect 39580 1912 39632 1921
rect 40316 1955 40368 1964
rect 40316 1921 40325 1955
rect 40325 1921 40359 1955
rect 40359 1921 40368 1955
rect 40316 1912 40368 1921
rect 41420 1912 41472 1964
rect 44916 1912 44968 1964
rect 30380 1844 30432 1896
rect 32220 1844 32272 1896
rect 34060 1844 34112 1896
rect 36820 1844 36872 1896
rect 39120 1844 39172 1896
rect 42340 1844 42392 1896
rect 43720 1844 43772 1896
rect 45928 1955 45980 1964
rect 45928 1921 45937 1955
rect 45937 1921 45971 1955
rect 45971 1921 45980 1955
rect 45928 1912 45980 1921
rect 46848 1955 46900 1964
rect 46848 1921 46857 1955
rect 46857 1921 46891 1955
rect 46891 1921 46900 1955
rect 46848 1912 46900 1921
rect 47032 1912 47084 1964
rect 46664 1887 46716 1896
rect 46664 1853 46673 1887
rect 46673 1853 46707 1887
rect 46707 1853 46716 1887
rect 46664 1844 46716 1853
rect 47860 1844 47912 1896
rect 22836 1751 22888 1760
rect 22836 1717 22845 1751
rect 22845 1717 22879 1751
rect 22879 1717 22888 1751
rect 22836 1708 22888 1717
rect 27804 1776 27856 1828
rect 28264 1776 28316 1828
rect 49424 2023 49476 2032
rect 49424 1989 49433 2023
rect 49433 1989 49467 2023
rect 49467 1989 49476 2023
rect 49424 1980 49476 1989
rect 51172 1980 51224 2032
rect 49608 1912 49660 1964
rect 49884 1912 49936 1964
rect 52460 1980 52512 2032
rect 52644 2023 52696 2032
rect 52644 1989 52653 2023
rect 52653 1989 52687 2023
rect 52687 1989 52696 2023
rect 52644 1980 52696 1989
rect 52276 1912 52328 1964
rect 50620 1844 50672 1896
rect 53196 1955 53248 1964
rect 53196 1921 53205 1955
rect 53205 1921 53239 1955
rect 53239 1921 53248 1955
rect 53196 1912 53248 1921
rect 53380 1844 53432 1896
rect 54944 1955 54996 1964
rect 54944 1921 54953 1955
rect 54953 1921 54987 1955
rect 54987 1921 54996 1955
rect 54944 1912 54996 1921
rect 55312 1912 55364 1964
rect 56048 1955 56100 1964
rect 56048 1921 56057 1955
rect 56057 1921 56091 1955
rect 56091 1921 56100 1955
rect 56048 1912 56100 1921
rect 57612 1955 57664 1964
rect 57612 1921 57621 1955
rect 57621 1921 57655 1955
rect 57655 1921 57664 1955
rect 57612 1912 57664 1921
rect 60464 1912 60516 1964
rect 61200 1955 61252 1964
rect 61200 1921 61209 1955
rect 61209 1921 61243 1955
rect 61243 1921 61252 1955
rect 61200 1912 61252 1921
rect 62488 1955 62540 1964
rect 62488 1921 62497 1955
rect 62497 1921 62531 1955
rect 62531 1921 62540 1955
rect 62488 1912 62540 1921
rect 56140 1844 56192 1896
rect 56968 1844 57020 1896
rect 58900 1844 58952 1896
rect 59544 1844 59596 1896
rect 62672 1844 62724 1896
rect 63040 1844 63092 1896
rect 64604 1955 64656 1964
rect 64604 1921 64613 1955
rect 64613 1921 64647 1955
rect 64647 1921 64656 1955
rect 64604 1912 64656 1921
rect 64788 1844 64840 1896
rect 24860 1708 24912 1760
rect 31392 1708 31444 1760
rect 40500 1751 40552 1760
rect 40500 1717 40509 1751
rect 40509 1717 40543 1751
rect 40543 1717 40552 1751
rect 40500 1708 40552 1717
rect 43260 1708 43312 1760
rect 46664 1708 46716 1760
rect 47308 1708 47360 1760
rect 47676 1751 47728 1760
rect 47676 1717 47685 1751
rect 47685 1717 47719 1751
rect 47719 1717 47728 1751
rect 47676 1708 47728 1717
rect 62396 1776 62448 1828
rect 63960 1776 64012 1828
rect 66812 1955 66864 1964
rect 66812 1921 66821 1955
rect 66821 1921 66855 1955
rect 66855 1921 66864 1955
rect 66812 1912 66864 1921
rect 68100 1955 68152 1964
rect 68100 1921 68109 1955
rect 68109 1921 68143 1955
rect 68143 1921 68152 1955
rect 68100 1912 68152 1921
rect 68284 1980 68336 2032
rect 72332 2048 72384 2100
rect 71136 2023 71188 2032
rect 71136 1989 71145 2023
rect 71145 1989 71179 2023
rect 71179 1989 71188 2023
rect 71136 1980 71188 1989
rect 73436 2023 73488 2032
rect 73436 1989 73445 2023
rect 73445 1989 73479 2023
rect 73479 1989 73488 2023
rect 73436 1980 73488 1989
rect 68652 1955 68704 1964
rect 68652 1921 68661 1955
rect 68661 1921 68695 1955
rect 68695 1921 68704 1955
rect 68652 1912 68704 1921
rect 70676 1955 70728 1964
rect 70676 1921 70685 1955
rect 70685 1921 70719 1955
rect 70719 1921 70728 1955
rect 70676 1912 70728 1921
rect 70860 1955 70912 1964
rect 70860 1921 70869 1955
rect 70869 1921 70903 1955
rect 70903 1921 70912 1955
rect 70860 1912 70912 1921
rect 71688 1912 71740 1964
rect 73712 1955 73764 1964
rect 73712 1921 73721 1955
rect 73721 1921 73755 1955
rect 73755 1921 73764 1955
rect 73712 1912 73764 1921
rect 68560 1844 68612 1896
rect 71320 1844 71372 1896
rect 70952 1776 71004 1828
rect 63868 1708 63920 1760
rect 67456 1751 67508 1760
rect 67456 1717 67465 1751
rect 67465 1717 67499 1751
rect 67499 1717 67508 1751
rect 67456 1708 67508 1717
rect 1858 1606 1910 1658
rect 1922 1606 1974 1658
rect 1986 1606 2038 1658
rect 2050 1606 2102 1658
rect 2114 1606 2166 1658
rect 11858 1606 11910 1658
rect 11922 1606 11974 1658
rect 11986 1606 12038 1658
rect 12050 1606 12102 1658
rect 12114 1606 12166 1658
rect 21858 1606 21910 1658
rect 21922 1606 21974 1658
rect 21986 1606 22038 1658
rect 22050 1606 22102 1658
rect 22114 1606 22166 1658
rect 31858 1606 31910 1658
rect 31922 1606 31974 1658
rect 31986 1606 32038 1658
rect 32050 1606 32102 1658
rect 32114 1606 32166 1658
rect 41858 1606 41910 1658
rect 41922 1606 41974 1658
rect 41986 1606 42038 1658
rect 42050 1606 42102 1658
rect 42114 1606 42166 1658
rect 51858 1606 51910 1658
rect 51922 1606 51974 1658
rect 51986 1606 52038 1658
rect 52050 1606 52102 1658
rect 52114 1606 52166 1658
rect 61858 1606 61910 1658
rect 61922 1606 61974 1658
rect 61986 1606 62038 1658
rect 62050 1606 62102 1658
rect 62114 1606 62166 1658
rect 71858 1606 71910 1658
rect 71922 1606 71974 1658
rect 71986 1606 72038 1658
rect 72050 1606 72102 1658
rect 72114 1606 72166 1658
rect 23572 1504 23624 1556
rect 33048 1504 33100 1556
rect 35532 1504 35584 1556
rect 41328 1504 41380 1556
rect 45560 1504 45612 1556
rect 46940 1504 46992 1556
rect 59728 1504 59780 1556
rect 20996 1343 21048 1352
rect 20996 1309 21005 1343
rect 21005 1309 21039 1343
rect 21039 1309 21048 1343
rect 20996 1300 21048 1309
rect 21732 1343 21784 1352
rect 21732 1309 21741 1343
rect 21741 1309 21775 1343
rect 21775 1309 21784 1343
rect 21732 1300 21784 1309
rect 22376 1368 22428 1420
rect 26148 1436 26200 1488
rect 30840 1436 30892 1488
rect 35624 1436 35676 1488
rect 65064 1504 65116 1556
rect 68468 1504 68520 1556
rect 73712 1504 73764 1556
rect 61660 1436 61712 1488
rect 22836 1411 22888 1420
rect 22836 1377 22845 1411
rect 22845 1377 22879 1411
rect 22879 1377 22888 1411
rect 22836 1368 22888 1377
rect 25136 1300 25188 1352
rect 25596 1343 25648 1352
rect 25596 1309 25605 1343
rect 25605 1309 25639 1343
rect 25639 1309 25648 1343
rect 25596 1300 25648 1309
rect 26424 1343 26476 1352
rect 26424 1309 26433 1343
rect 26433 1309 26467 1343
rect 26467 1309 26476 1343
rect 26424 1300 26476 1309
rect 26700 1343 26752 1352
rect 26700 1309 26709 1343
rect 26709 1309 26743 1343
rect 26743 1309 26752 1343
rect 26700 1300 26752 1309
rect 27160 1343 27212 1352
rect 27160 1309 27169 1343
rect 27169 1309 27203 1343
rect 27203 1309 27212 1343
rect 27160 1300 27212 1309
rect 20812 1207 20864 1216
rect 20812 1173 20821 1207
rect 20821 1173 20855 1207
rect 20855 1173 20864 1207
rect 20812 1164 20864 1173
rect 21548 1207 21600 1216
rect 21548 1173 21557 1207
rect 21557 1173 21591 1207
rect 21591 1173 21600 1207
rect 21548 1164 21600 1173
rect 22284 1164 22336 1216
rect 22652 1207 22704 1216
rect 22652 1173 22661 1207
rect 22661 1173 22695 1207
rect 22695 1173 22704 1207
rect 22652 1164 22704 1173
rect 23388 1207 23440 1216
rect 23388 1173 23397 1207
rect 23397 1173 23431 1207
rect 23431 1173 23440 1207
rect 23388 1164 23440 1173
rect 23940 1232 23992 1284
rect 28540 1232 28592 1284
rect 29276 1343 29328 1352
rect 29276 1309 29285 1343
rect 29285 1309 29319 1343
rect 29319 1309 29328 1343
rect 29276 1300 29328 1309
rect 30748 1232 30800 1284
rect 26884 1164 26936 1216
rect 30472 1164 30524 1216
rect 31576 1300 31628 1352
rect 32956 1343 33008 1352
rect 32956 1309 32965 1343
rect 32965 1309 32999 1343
rect 32999 1309 33008 1343
rect 32956 1300 33008 1309
rect 38660 1368 38712 1420
rect 33508 1164 33560 1216
rect 33968 1275 34020 1284
rect 33968 1241 33977 1275
rect 33977 1241 34011 1275
rect 34011 1241 34020 1275
rect 33968 1232 34020 1241
rect 35072 1232 35124 1284
rect 35440 1232 35492 1284
rect 36544 1232 36596 1284
rect 36912 1343 36964 1352
rect 36912 1309 36921 1343
rect 36921 1309 36955 1343
rect 36955 1309 36964 1343
rect 36912 1300 36964 1309
rect 37280 1232 37332 1284
rect 38200 1232 38252 1284
rect 39396 1343 39448 1352
rect 39396 1309 39405 1343
rect 39405 1309 39439 1343
rect 39439 1309 39448 1343
rect 39396 1300 39448 1309
rect 40500 1300 40552 1352
rect 41144 1343 41196 1352
rect 41144 1309 41153 1343
rect 41153 1309 41187 1343
rect 41187 1309 41196 1343
rect 41144 1300 41196 1309
rect 42800 1368 42852 1420
rect 43996 1300 44048 1352
rect 44824 1300 44876 1352
rect 46388 1343 46440 1352
rect 46388 1309 46397 1343
rect 46397 1309 46431 1343
rect 46431 1309 46440 1343
rect 46388 1300 46440 1309
rect 48504 1368 48556 1420
rect 49056 1300 49108 1352
rect 49332 1300 49384 1352
rect 51448 1343 51500 1352
rect 51448 1309 51457 1343
rect 51457 1309 51491 1343
rect 51491 1309 51500 1343
rect 51448 1300 51500 1309
rect 55864 1368 55916 1420
rect 65156 1436 65208 1488
rect 64972 1411 65024 1420
rect 64972 1377 64981 1411
rect 64981 1377 65015 1411
rect 65015 1377 65024 1411
rect 64972 1368 65024 1377
rect 67180 1368 67232 1420
rect 69940 1368 69992 1420
rect 74632 1411 74684 1420
rect 74632 1377 74641 1411
rect 74641 1377 74675 1411
rect 74675 1377 74684 1411
rect 74632 1368 74684 1377
rect 51632 1300 51684 1352
rect 54024 1343 54076 1352
rect 54024 1309 54033 1343
rect 54033 1309 54067 1343
rect 54067 1309 54076 1343
rect 54024 1300 54076 1309
rect 39580 1232 39632 1284
rect 40132 1232 40184 1284
rect 41328 1232 41380 1284
rect 45100 1232 45152 1284
rect 46480 1232 46532 1284
rect 48320 1232 48372 1284
rect 49240 1232 49292 1284
rect 41052 1164 41104 1216
rect 50160 1164 50212 1216
rect 52368 1232 52420 1284
rect 54760 1232 54812 1284
rect 53932 1164 53984 1216
rect 56692 1343 56744 1352
rect 56692 1309 56701 1343
rect 56701 1309 56735 1343
rect 56735 1309 56744 1343
rect 56692 1300 56744 1309
rect 57244 1343 57296 1352
rect 57244 1309 57253 1343
rect 57253 1309 57287 1343
rect 57287 1309 57296 1343
rect 57244 1300 57296 1309
rect 59084 1343 59136 1352
rect 59084 1309 59093 1343
rect 59093 1309 59127 1343
rect 59127 1309 59136 1343
rect 59084 1300 59136 1309
rect 59268 1343 59320 1352
rect 59268 1309 59277 1343
rect 59277 1309 59311 1343
rect 59311 1309 59320 1343
rect 59268 1300 59320 1309
rect 59452 1300 59504 1352
rect 62304 1300 62356 1352
rect 62396 1343 62448 1352
rect 62396 1309 62405 1343
rect 62405 1309 62439 1343
rect 62439 1309 62448 1343
rect 62396 1300 62448 1309
rect 63132 1343 63184 1352
rect 63132 1309 63141 1343
rect 63141 1309 63175 1343
rect 63175 1309 63184 1343
rect 63132 1300 63184 1309
rect 63408 1300 63460 1352
rect 65892 1343 65944 1352
rect 65892 1309 65901 1343
rect 65901 1309 65935 1343
rect 65935 1309 65944 1343
rect 65892 1300 65944 1309
rect 67456 1343 67508 1352
rect 67456 1309 67465 1343
rect 67465 1309 67499 1343
rect 67499 1309 67508 1343
rect 67456 1300 67508 1309
rect 68192 1343 68244 1352
rect 68192 1309 68201 1343
rect 68201 1309 68235 1343
rect 68235 1309 68244 1343
rect 68192 1300 68244 1309
rect 69388 1300 69440 1352
rect 69756 1300 69808 1352
rect 70768 1343 70820 1352
rect 70768 1309 70777 1343
rect 70777 1309 70811 1343
rect 70811 1309 70820 1343
rect 70768 1300 70820 1309
rect 72240 1300 72292 1352
rect 72700 1343 72752 1352
rect 72700 1309 72709 1343
rect 72709 1309 72743 1343
rect 72743 1309 72752 1343
rect 72700 1300 72752 1309
rect 73252 1343 73304 1352
rect 73252 1309 73261 1343
rect 73261 1309 73295 1343
rect 73295 1309 73304 1343
rect 73252 1300 73304 1309
rect 57520 1232 57572 1284
rect 60280 1232 60332 1284
rect 61660 1232 61712 1284
rect 65800 1232 65852 1284
rect 70860 1232 70912 1284
rect 63684 1164 63736 1216
rect 4210 1062 4262 1114
rect 4274 1062 4326 1114
rect 4338 1062 4390 1114
rect 4402 1062 4454 1114
rect 4466 1062 4518 1114
rect 14210 1062 14262 1114
rect 14274 1062 14326 1114
rect 14338 1062 14390 1114
rect 14402 1062 14454 1114
rect 14466 1062 14518 1114
rect 24210 1062 24262 1114
rect 24274 1062 24326 1114
rect 24338 1062 24390 1114
rect 24402 1062 24454 1114
rect 24466 1062 24518 1114
rect 34210 1062 34262 1114
rect 34274 1062 34326 1114
rect 34338 1062 34390 1114
rect 34402 1062 34454 1114
rect 34466 1062 34518 1114
rect 44210 1062 44262 1114
rect 44274 1062 44326 1114
rect 44338 1062 44390 1114
rect 44402 1062 44454 1114
rect 44466 1062 44518 1114
rect 54210 1062 54262 1114
rect 54274 1062 54326 1114
rect 54338 1062 54390 1114
rect 54402 1062 54454 1114
rect 54466 1062 54518 1114
rect 64210 1062 64262 1114
rect 64274 1062 64326 1114
rect 64338 1062 64390 1114
rect 64402 1062 64454 1114
rect 64466 1062 64518 1114
rect 74210 1062 74262 1114
rect 74274 1062 74326 1114
rect 74338 1062 74390 1114
rect 74402 1062 74454 1114
rect 74466 1062 74518 1114
rect 21732 960 21784 1012
rect 23296 960 23348 1012
rect 23388 960 23440 1012
rect 26516 960 26568 1012
rect 30472 960 30524 1012
rect 33876 960 33928 1012
rect 36544 960 36596 1012
rect 39764 960 39816 1012
rect 41144 960 41196 1012
rect 65984 960 66036 1012
rect 20812 892 20864 944
rect 23664 892 23716 944
rect 29000 892 29052 944
rect 33968 892 34020 944
rect 40408 892 40460 944
rect 49056 892 49108 944
rect 72608 892 72660 944
rect 22376 824 22428 876
rect 26056 824 26108 876
rect 21548 756 21600 808
rect 25044 756 25096 808
rect 25136 756 25188 808
rect 43996 824 44048 876
rect 65432 824 65484 876
rect 29276 756 29328 808
rect 64052 756 64104 808
rect 22652 688 22704 740
rect 28356 688 28408 740
rect 46388 688 46440 740
rect 70492 688 70544 740
rect 36912 620 36964 672
rect 65248 620 65300 672
rect 39396 552 39448 604
rect 64972 552 65024 604
rect 54024 484 54076 536
rect 63776 484 63828 536
rect 63132 348 63184 400
rect 72792 348 72844 400
rect 51448 280 51500 332
rect 65616 280 65668 332
<< metal2 >>
rect 71836 85434 72188 86000
rect 71836 85382 71858 85434
rect 71910 85382 71922 85434
rect 71974 85382 71986 85434
rect 72038 85382 72050 85434
rect 72102 85382 72114 85434
rect 72166 85382 72188 85434
rect 2020 84588 2124 84616
rect 2020 84532 2044 84588
rect 2100 84532 2124 84588
rect 2020 84508 2124 84532
rect 2020 84452 2044 84508
rect 2100 84452 2124 84508
rect 2020 84428 2124 84452
rect 2020 84372 2044 84428
rect 2100 84372 2124 84428
rect 2020 84348 2124 84372
rect 2020 84292 2044 84348
rect 2100 84292 2124 84348
rect 2020 84264 2124 84292
rect 5521 84588 5615 84616
rect 5521 84532 5540 84588
rect 5596 84532 5615 84588
rect 5521 84508 5615 84532
rect 5521 84452 5540 84508
rect 5596 84452 5615 84508
rect 5521 84428 5615 84452
rect 5521 84372 5540 84428
rect 5596 84372 5615 84428
rect 5521 84348 5615 84372
rect 5521 84292 5540 84348
rect 5596 84292 5615 84348
rect 5521 84264 5615 84292
rect 8411 84588 8505 84616
rect 8411 84532 8430 84588
rect 8486 84532 8505 84588
rect 8411 84508 8505 84532
rect 8411 84452 8430 84508
rect 8486 84452 8505 84508
rect 8411 84428 8505 84452
rect 8411 84372 8430 84428
rect 8486 84372 8505 84428
rect 8411 84348 8505 84372
rect 8411 84292 8430 84348
rect 8486 84292 8505 84348
rect 8411 84264 8505 84292
rect 11301 84588 11395 84616
rect 11301 84532 11320 84588
rect 11376 84532 11395 84588
rect 11301 84508 11395 84532
rect 11301 84452 11320 84508
rect 11376 84452 11395 84508
rect 11301 84428 11395 84452
rect 11301 84372 11320 84428
rect 11376 84372 11395 84428
rect 11301 84348 11395 84372
rect 11301 84292 11320 84348
rect 11376 84292 11395 84348
rect 11301 84264 11395 84292
rect 14191 84588 14285 84616
rect 14191 84532 14210 84588
rect 14266 84532 14285 84588
rect 14191 84508 14285 84532
rect 14191 84452 14210 84508
rect 14266 84452 14285 84508
rect 14191 84428 14285 84452
rect 14191 84372 14210 84428
rect 14266 84372 14285 84428
rect 14191 84348 14285 84372
rect 14191 84292 14210 84348
rect 14266 84292 14285 84348
rect 14191 84264 14285 84292
rect 17081 84588 17175 84616
rect 17081 84532 17100 84588
rect 17156 84532 17175 84588
rect 17081 84508 17175 84532
rect 17081 84452 17100 84508
rect 17156 84452 17175 84508
rect 17081 84428 17175 84452
rect 17081 84372 17100 84428
rect 17156 84372 17175 84428
rect 17081 84348 17175 84372
rect 17081 84292 17100 84348
rect 17156 84292 17175 84348
rect 17081 84264 17175 84292
rect 19971 84588 20065 84616
rect 19971 84532 19990 84588
rect 20046 84532 20065 84588
rect 19971 84508 20065 84532
rect 19971 84452 19990 84508
rect 20046 84452 20065 84508
rect 19971 84428 20065 84452
rect 19971 84372 19990 84428
rect 20046 84372 20065 84428
rect 19971 84348 20065 84372
rect 19971 84292 19990 84348
rect 20046 84292 20065 84348
rect 19971 84264 20065 84292
rect 22861 84588 22955 84616
rect 22861 84532 22880 84588
rect 22936 84532 22955 84588
rect 22861 84508 22955 84532
rect 22861 84452 22880 84508
rect 22936 84452 22955 84508
rect 22861 84428 22955 84452
rect 22861 84372 22880 84428
rect 22936 84372 22955 84428
rect 22861 84348 22955 84372
rect 22861 84292 22880 84348
rect 22936 84292 22955 84348
rect 22861 84264 22955 84292
rect 25751 84588 25845 84616
rect 25751 84532 25770 84588
rect 25826 84532 25845 84588
rect 25751 84508 25845 84532
rect 25751 84452 25770 84508
rect 25826 84452 25845 84508
rect 25751 84428 25845 84452
rect 25751 84372 25770 84428
rect 25826 84372 25845 84428
rect 25751 84348 25845 84372
rect 25751 84292 25770 84348
rect 25826 84292 25845 84348
rect 25751 84264 25845 84292
rect 28641 84588 28735 84616
rect 28641 84532 28660 84588
rect 28716 84532 28735 84588
rect 28641 84508 28735 84532
rect 28641 84452 28660 84508
rect 28716 84452 28735 84508
rect 28641 84428 28735 84452
rect 28641 84372 28660 84428
rect 28716 84372 28735 84428
rect 28641 84348 28735 84372
rect 28641 84292 28660 84348
rect 28716 84292 28735 84348
rect 28641 84264 28735 84292
rect 31531 84588 31625 84616
rect 31531 84532 31550 84588
rect 31606 84532 31625 84588
rect 31531 84508 31625 84532
rect 31531 84452 31550 84508
rect 31606 84452 31625 84508
rect 31531 84428 31625 84452
rect 31531 84372 31550 84428
rect 31606 84372 31625 84428
rect 31531 84348 31625 84372
rect 31531 84292 31550 84348
rect 31606 84292 31625 84348
rect 31531 84264 31625 84292
rect 34421 84588 34515 84616
rect 34421 84532 34440 84588
rect 34496 84532 34515 84588
rect 34421 84508 34515 84532
rect 34421 84452 34440 84508
rect 34496 84452 34515 84508
rect 34421 84428 34515 84452
rect 34421 84372 34440 84428
rect 34496 84372 34515 84428
rect 34421 84348 34515 84372
rect 34421 84292 34440 84348
rect 34496 84292 34515 84348
rect 34421 84264 34515 84292
rect 37311 84588 37405 84616
rect 37311 84532 37330 84588
rect 37386 84532 37405 84588
rect 37311 84508 37405 84532
rect 37311 84452 37330 84508
rect 37386 84452 37405 84508
rect 37311 84428 37405 84452
rect 37311 84372 37330 84428
rect 37386 84372 37405 84428
rect 37311 84348 37405 84372
rect 37311 84292 37330 84348
rect 37386 84292 37405 84348
rect 37311 84264 37405 84292
rect 40201 84588 40295 84616
rect 40201 84532 40220 84588
rect 40276 84532 40295 84588
rect 40201 84508 40295 84532
rect 40201 84452 40220 84508
rect 40276 84452 40295 84508
rect 40201 84428 40295 84452
rect 40201 84372 40220 84428
rect 40276 84372 40295 84428
rect 40201 84348 40295 84372
rect 40201 84292 40220 84348
rect 40276 84292 40295 84348
rect 40201 84264 40295 84292
rect 43091 84588 43185 84616
rect 43091 84532 43110 84588
rect 43166 84532 43185 84588
rect 43091 84508 43185 84532
rect 43091 84452 43110 84508
rect 43166 84452 43185 84508
rect 43091 84428 43185 84452
rect 43091 84372 43110 84428
rect 43166 84372 43185 84428
rect 43091 84348 43185 84372
rect 43091 84292 43110 84348
rect 43166 84292 43185 84348
rect 43091 84264 43185 84292
rect 45981 84588 46075 84616
rect 45981 84532 46000 84588
rect 46056 84532 46075 84588
rect 45981 84508 46075 84532
rect 45981 84452 46000 84508
rect 46056 84452 46075 84508
rect 45981 84428 46075 84452
rect 45981 84372 46000 84428
rect 46056 84372 46075 84428
rect 45981 84348 46075 84372
rect 45981 84292 46000 84348
rect 46056 84292 46075 84348
rect 45981 84264 46075 84292
rect 48989 84588 49083 84616
rect 48989 84532 49008 84588
rect 49064 84532 49083 84588
rect 48989 84508 49083 84532
rect 48989 84452 49008 84508
rect 49064 84452 49083 84508
rect 48989 84428 49083 84452
rect 48989 84372 49008 84428
rect 49064 84372 49083 84428
rect 48989 84348 49083 84372
rect 48989 84292 49008 84348
rect 49064 84292 49083 84348
rect 48989 84264 49083 84292
rect 52210 84588 52320 84616
rect 52210 84532 52237 84588
rect 52293 84532 52320 84588
rect 52210 84508 52320 84532
rect 52210 84452 52237 84508
rect 52293 84452 52320 84508
rect 52210 84428 52320 84452
rect 52210 84372 52237 84428
rect 52293 84372 52320 84428
rect 52210 84348 52320 84372
rect 52210 84292 52237 84348
rect 52293 84292 52320 84348
rect 52210 84264 52320 84292
rect 53602 84588 53730 84616
rect 53602 84532 53638 84588
rect 53694 84532 53730 84588
rect 53602 84508 53730 84532
rect 53602 84452 53638 84508
rect 53694 84452 53730 84508
rect 53602 84428 53730 84452
rect 53602 84372 53638 84428
rect 53694 84372 53730 84428
rect 53602 84348 53730 84372
rect 53602 84292 53638 84348
rect 53694 84292 53730 84348
rect 53602 84264 53730 84292
rect 53770 84588 53898 84616
rect 53770 84532 53806 84588
rect 53862 84532 53898 84588
rect 53770 84508 53898 84532
rect 53770 84452 53806 84508
rect 53862 84452 53898 84508
rect 53770 84428 53898 84452
rect 53770 84372 53806 84428
rect 53862 84372 53898 84428
rect 53770 84348 53898 84372
rect 53770 84292 53806 84348
rect 53862 84292 53898 84348
rect 53770 84264 53898 84292
rect 54514 84588 54642 84616
rect 54514 84532 54550 84588
rect 54606 84532 54642 84588
rect 54514 84508 54642 84532
rect 54514 84452 54550 84508
rect 54606 84452 54642 84508
rect 54514 84428 54642 84452
rect 54514 84372 54550 84428
rect 54606 84372 54642 84428
rect 54514 84348 54642 84372
rect 54514 84292 54550 84348
rect 54606 84292 54642 84348
rect 54514 84264 54642 84292
rect 54910 84588 55026 84616
rect 54910 84532 54940 84588
rect 54996 84532 55026 84588
rect 54910 84508 55026 84532
rect 54910 84452 54940 84508
rect 54996 84452 55026 84508
rect 54910 84428 55026 84452
rect 54910 84372 54940 84428
rect 54996 84372 55026 84428
rect 54910 84348 55026 84372
rect 54910 84292 54940 84348
rect 54996 84292 55026 84348
rect 54910 84264 55026 84292
rect 55620 84588 55748 84616
rect 55620 84532 55656 84588
rect 55712 84532 55748 84588
rect 55620 84508 55748 84532
rect 55620 84452 55656 84508
rect 55712 84452 55748 84508
rect 55620 84428 55748 84452
rect 55620 84372 55656 84428
rect 55712 84372 55748 84428
rect 55620 84348 55748 84372
rect 55620 84292 55656 84348
rect 55712 84292 55748 84348
rect 55620 84264 55748 84292
rect 56198 84588 56326 84616
rect 56198 84532 56234 84588
rect 56290 84532 56326 84588
rect 56198 84508 56326 84532
rect 56198 84452 56234 84508
rect 56290 84452 56326 84508
rect 56198 84428 56326 84452
rect 56198 84372 56234 84428
rect 56290 84372 56326 84428
rect 56198 84348 56326 84372
rect 56198 84292 56234 84348
rect 56290 84292 56326 84348
rect 56198 84264 56326 84292
rect 56649 84588 56765 84616
rect 56649 84532 56679 84588
rect 56735 84532 56765 84588
rect 56649 84508 56765 84532
rect 56649 84452 56679 84508
rect 56735 84452 56765 84508
rect 56649 84428 56765 84452
rect 56649 84372 56679 84428
rect 56735 84372 56765 84428
rect 56649 84348 56765 84372
rect 56649 84292 56679 84348
rect 56735 84292 56765 84348
rect 56649 84264 56765 84292
rect 56953 84588 57069 84616
rect 56953 84532 56983 84588
rect 57039 84532 57069 84588
rect 56953 84508 57069 84532
rect 56953 84452 56983 84508
rect 57039 84452 57069 84508
rect 56953 84428 57069 84452
rect 56953 84372 56983 84428
rect 57039 84372 57069 84428
rect 56953 84348 57069 84372
rect 56953 84292 56983 84348
rect 57039 84292 57069 84348
rect 56953 84264 57069 84292
rect 57795 84588 57911 84616
rect 57795 84532 57825 84588
rect 57881 84532 57911 84588
rect 57795 84508 57911 84532
rect 57795 84452 57825 84508
rect 57881 84452 57911 84508
rect 57795 84428 57911 84452
rect 57795 84372 57825 84428
rect 57881 84372 57911 84428
rect 57795 84348 57911 84372
rect 57795 84292 57825 84348
rect 57881 84292 57911 84348
rect 57795 84264 57911 84292
rect 58461 84588 58525 84616
rect 58461 84532 58465 84588
rect 58521 84532 58525 84588
rect 58461 84508 58525 84532
rect 58461 84452 58465 84508
rect 58521 84452 58525 84508
rect 58461 84428 58525 84452
rect 58461 84372 58465 84428
rect 58521 84372 58525 84428
rect 58461 84348 58525 84372
rect 58461 84292 58465 84348
rect 58521 84292 58525 84348
rect 58461 84264 58525 84292
rect 59018 84588 59134 84616
rect 59018 84532 59048 84588
rect 59104 84532 59134 84588
rect 59018 84508 59134 84532
rect 59018 84452 59048 84508
rect 59104 84452 59134 84508
rect 59018 84428 59134 84452
rect 59018 84372 59048 84428
rect 59104 84372 59134 84428
rect 59018 84348 59134 84372
rect 59018 84292 59048 84348
rect 59104 84292 59134 84348
rect 59018 84264 59134 84292
rect 60296 84588 60412 84616
rect 60296 84532 60326 84588
rect 60382 84532 60412 84588
rect 60296 84508 60412 84532
rect 60296 84452 60326 84508
rect 60382 84452 60412 84508
rect 60296 84428 60412 84452
rect 60296 84372 60326 84428
rect 60382 84372 60412 84428
rect 60296 84348 60412 84372
rect 60296 84292 60326 84348
rect 60382 84292 60412 84348
rect 60296 84264 60412 84292
rect 60454 84588 60570 84616
rect 60454 84532 60484 84588
rect 60540 84532 60570 84588
rect 60454 84508 60570 84532
rect 60454 84452 60484 84508
rect 60540 84452 60570 84508
rect 60454 84428 60570 84452
rect 60454 84372 60484 84428
rect 60540 84372 60570 84428
rect 60454 84348 60570 84372
rect 60454 84292 60484 84348
rect 60540 84292 60570 84348
rect 60454 84264 60570 84292
rect 62509 84588 62683 84616
rect 62509 84532 62528 84588
rect 62584 84532 62608 84588
rect 62664 84532 62683 84588
rect 62509 84508 62683 84532
rect 62509 84452 62528 84508
rect 62584 84452 62608 84508
rect 62664 84452 62683 84508
rect 62509 84428 62683 84452
rect 62509 84372 62528 84428
rect 62584 84372 62608 84428
rect 62664 84372 62683 84428
rect 62509 84348 62683 84372
rect 62509 84292 62528 84348
rect 62584 84292 62608 84348
rect 62664 84292 62683 84348
rect 62509 84264 62683 84292
rect 71836 84346 72188 85382
rect 71836 84294 71858 84346
rect 71910 84294 71922 84346
rect 71974 84294 71986 84346
rect 72038 84294 72050 84346
rect 72102 84294 72114 84346
rect 72166 84294 72188 84346
rect 64880 84244 64932 84250
rect 64880 84186 64932 84192
rect 2152 82236 2352 82264
rect 2152 82180 2184 82236
rect 2240 82180 2264 82236
rect 2320 82180 2352 82236
rect 2152 82156 2352 82180
rect 2152 82100 2184 82156
rect 2240 82100 2264 82156
rect 2320 82100 2352 82156
rect 2152 82076 2352 82100
rect 2152 82020 2184 82076
rect 2240 82020 2264 82076
rect 2320 82020 2352 82076
rect 2152 81996 2352 82020
rect 2152 81940 2184 81996
rect 2240 81940 2264 81996
rect 2320 81940 2352 81996
rect 2152 81912 2352 81940
rect 5374 82236 5468 82264
rect 5374 82180 5393 82236
rect 5449 82180 5468 82236
rect 5374 82156 5468 82180
rect 5374 82100 5393 82156
rect 5449 82100 5468 82156
rect 5374 82076 5468 82100
rect 5374 82020 5393 82076
rect 5449 82020 5468 82076
rect 5374 81996 5468 82020
rect 5374 81940 5393 81996
rect 5449 81940 5468 81996
rect 5374 81912 5468 81940
rect 8264 82236 8358 82264
rect 8264 82180 8283 82236
rect 8339 82180 8358 82236
rect 8264 82156 8358 82180
rect 8264 82100 8283 82156
rect 8339 82100 8358 82156
rect 8264 82076 8358 82100
rect 8264 82020 8283 82076
rect 8339 82020 8358 82076
rect 8264 81996 8358 82020
rect 8264 81940 8283 81996
rect 8339 81940 8358 81996
rect 8264 81912 8358 81940
rect 11154 82236 11248 82264
rect 11154 82180 11173 82236
rect 11229 82180 11248 82236
rect 11154 82156 11248 82180
rect 11154 82100 11173 82156
rect 11229 82100 11248 82156
rect 11154 82076 11248 82100
rect 11154 82020 11173 82076
rect 11229 82020 11248 82076
rect 11154 81996 11248 82020
rect 11154 81940 11173 81996
rect 11229 81940 11248 81996
rect 11154 81912 11248 81940
rect 14044 82236 14138 82264
rect 14044 82180 14063 82236
rect 14119 82180 14138 82236
rect 14044 82156 14138 82180
rect 14044 82100 14063 82156
rect 14119 82100 14138 82156
rect 14044 82076 14138 82100
rect 14044 82020 14063 82076
rect 14119 82020 14138 82076
rect 14044 81996 14138 82020
rect 14044 81940 14063 81996
rect 14119 81940 14138 81996
rect 14044 81912 14138 81940
rect 16934 82236 17028 82264
rect 16934 82180 16953 82236
rect 17009 82180 17028 82236
rect 16934 82156 17028 82180
rect 16934 82100 16953 82156
rect 17009 82100 17028 82156
rect 16934 82076 17028 82100
rect 16934 82020 16953 82076
rect 17009 82020 17028 82076
rect 16934 81996 17028 82020
rect 16934 81940 16953 81996
rect 17009 81940 17028 81996
rect 16934 81912 17028 81940
rect 19824 82236 19918 82264
rect 19824 82180 19843 82236
rect 19899 82180 19918 82236
rect 19824 82156 19918 82180
rect 19824 82100 19843 82156
rect 19899 82100 19918 82156
rect 19824 82076 19918 82100
rect 19824 82020 19843 82076
rect 19899 82020 19918 82076
rect 19824 81996 19918 82020
rect 19824 81940 19843 81996
rect 19899 81940 19918 81996
rect 19824 81912 19918 81940
rect 22714 82236 22808 82264
rect 22714 82180 22733 82236
rect 22789 82180 22808 82236
rect 22714 82156 22808 82180
rect 22714 82100 22733 82156
rect 22789 82100 22808 82156
rect 22714 82076 22808 82100
rect 22714 82020 22733 82076
rect 22789 82020 22808 82076
rect 22714 81996 22808 82020
rect 22714 81940 22733 81996
rect 22789 81940 22808 81996
rect 22714 81912 22808 81940
rect 25604 82236 25698 82264
rect 25604 82180 25623 82236
rect 25679 82180 25698 82236
rect 25604 82156 25698 82180
rect 25604 82100 25623 82156
rect 25679 82100 25698 82156
rect 25604 82076 25698 82100
rect 25604 82020 25623 82076
rect 25679 82020 25698 82076
rect 25604 81996 25698 82020
rect 25604 81940 25623 81996
rect 25679 81940 25698 81996
rect 25604 81912 25698 81940
rect 28494 82236 28588 82264
rect 28494 82180 28513 82236
rect 28569 82180 28588 82236
rect 28494 82156 28588 82180
rect 28494 82100 28513 82156
rect 28569 82100 28588 82156
rect 28494 82076 28588 82100
rect 28494 82020 28513 82076
rect 28569 82020 28588 82076
rect 28494 81996 28588 82020
rect 28494 81940 28513 81996
rect 28569 81940 28588 81996
rect 28494 81912 28588 81940
rect 31384 82236 31478 82264
rect 31384 82180 31403 82236
rect 31459 82180 31478 82236
rect 31384 82156 31478 82180
rect 31384 82100 31403 82156
rect 31459 82100 31478 82156
rect 31384 82076 31478 82100
rect 31384 82020 31403 82076
rect 31459 82020 31478 82076
rect 31384 81996 31478 82020
rect 31384 81940 31403 81996
rect 31459 81940 31478 81996
rect 31384 81912 31478 81940
rect 34274 82236 34368 82264
rect 34274 82180 34293 82236
rect 34349 82180 34368 82236
rect 34274 82156 34368 82180
rect 34274 82100 34293 82156
rect 34349 82100 34368 82156
rect 34274 82076 34368 82100
rect 34274 82020 34293 82076
rect 34349 82020 34368 82076
rect 34274 81996 34368 82020
rect 34274 81940 34293 81996
rect 34349 81940 34368 81996
rect 34274 81912 34368 81940
rect 37164 82236 37258 82264
rect 37164 82180 37183 82236
rect 37239 82180 37258 82236
rect 37164 82156 37258 82180
rect 37164 82100 37183 82156
rect 37239 82100 37258 82156
rect 37164 82076 37258 82100
rect 37164 82020 37183 82076
rect 37239 82020 37258 82076
rect 37164 81996 37258 82020
rect 37164 81940 37183 81996
rect 37239 81940 37258 81996
rect 37164 81912 37258 81940
rect 40054 82236 40148 82264
rect 40054 82180 40073 82236
rect 40129 82180 40148 82236
rect 40054 82156 40148 82180
rect 40054 82100 40073 82156
rect 40129 82100 40148 82156
rect 40054 82076 40148 82100
rect 40054 82020 40073 82076
rect 40129 82020 40148 82076
rect 40054 81996 40148 82020
rect 40054 81940 40073 81996
rect 40129 81940 40148 81996
rect 40054 81912 40148 81940
rect 42944 82236 43038 82264
rect 42944 82180 42963 82236
rect 43019 82180 43038 82236
rect 42944 82156 43038 82180
rect 42944 82100 42963 82156
rect 43019 82100 43038 82156
rect 42944 82076 43038 82100
rect 42944 82020 42963 82076
rect 43019 82020 43038 82076
rect 42944 81996 43038 82020
rect 42944 81940 42963 81996
rect 43019 81940 43038 81996
rect 42944 81912 43038 81940
rect 45834 82236 45928 82264
rect 45834 82180 45853 82236
rect 45909 82180 45928 82236
rect 45834 82156 45928 82180
rect 45834 82100 45853 82156
rect 45909 82100 45928 82156
rect 45834 82076 45928 82100
rect 45834 82020 45853 82076
rect 45909 82020 45928 82076
rect 45834 81996 45928 82020
rect 45834 81940 45853 81996
rect 45909 81940 45928 81996
rect 45834 81912 45928 81940
rect 48781 82236 48875 82264
rect 48781 82180 48800 82236
rect 48856 82180 48875 82236
rect 48781 82156 48875 82180
rect 48781 82100 48800 82156
rect 48856 82100 48875 82156
rect 48781 82076 48875 82100
rect 48781 82020 48800 82076
rect 48856 82020 48875 82076
rect 48781 81996 48875 82020
rect 48781 81940 48800 81996
rect 48856 81940 48875 81996
rect 48781 81912 48875 81940
rect 49630 82236 49830 82264
rect 49630 82180 49662 82236
rect 49718 82180 49742 82236
rect 49798 82180 49830 82236
rect 49630 82156 49830 82180
rect 49630 82100 49662 82156
rect 49718 82100 49742 82156
rect 49798 82100 49830 82156
rect 49630 82076 49830 82100
rect 49630 82020 49662 82076
rect 49718 82020 49742 82076
rect 49798 82020 49830 82076
rect 49630 81996 49830 82020
rect 49630 81940 49662 81996
rect 49718 81940 49742 81996
rect 49798 81940 49830 81996
rect 49630 81912 49830 81940
rect 52920 82236 53048 82264
rect 52920 82180 52956 82236
rect 53012 82180 53048 82236
rect 52920 82156 53048 82180
rect 52920 82100 52956 82156
rect 53012 82100 53048 82156
rect 52920 82076 53048 82100
rect 52920 82020 52956 82076
rect 53012 82020 53048 82076
rect 52920 81996 53048 82020
rect 52920 81940 52956 81996
rect 53012 81940 53048 81996
rect 52920 81912 53048 81940
rect 53078 82236 53206 82264
rect 53078 82180 53114 82236
rect 53170 82180 53206 82236
rect 53078 82156 53206 82180
rect 53078 82100 53114 82156
rect 53170 82100 53206 82156
rect 53078 82076 53206 82100
rect 53078 82020 53114 82076
rect 53170 82020 53206 82076
rect 53078 81996 53206 82020
rect 53078 81940 53114 81996
rect 53170 81940 53206 81996
rect 53078 81912 53206 81940
rect 53434 82236 53562 82264
rect 53434 82180 53470 82236
rect 53526 82180 53562 82236
rect 53434 82156 53562 82180
rect 53434 82100 53470 82156
rect 53526 82100 53562 82156
rect 53434 82076 53562 82100
rect 53434 82020 53470 82076
rect 53526 82020 53562 82076
rect 53434 81996 53562 82020
rect 53434 81940 53470 81996
rect 53526 81940 53562 81996
rect 53434 81912 53562 81940
rect 54752 82236 54880 82264
rect 54752 82180 54788 82236
rect 54844 82180 54880 82236
rect 54752 82156 54880 82180
rect 54752 82100 54788 82156
rect 54844 82100 54880 82156
rect 54752 82076 54880 82100
rect 54752 82020 54788 82076
rect 54844 82020 54880 82076
rect 54752 81996 54880 82020
rect 54752 81940 54788 81996
rect 54844 81940 54880 81996
rect 54752 81912 54880 81940
rect 55345 82236 55473 82264
rect 55345 82180 55381 82236
rect 55437 82180 55473 82236
rect 55345 82156 55473 82180
rect 55345 82100 55381 82156
rect 55437 82100 55473 82156
rect 55345 82076 55473 82100
rect 55345 82020 55381 82076
rect 55437 82020 55473 82076
rect 55345 81996 55473 82020
rect 55345 81940 55381 81996
rect 55437 81940 55473 81996
rect 55345 81912 55473 81940
rect 56491 82236 56619 82264
rect 56491 82180 56527 82236
rect 56583 82180 56619 82236
rect 56491 82156 56619 82180
rect 56491 82100 56527 82156
rect 56583 82100 56619 82156
rect 56491 82076 56619 82100
rect 56491 82020 56527 82076
rect 56583 82020 56619 82076
rect 56491 81996 56619 82020
rect 56491 81940 56527 81996
rect 56583 81940 56619 81996
rect 56491 81912 56619 81940
rect 57941 82236 58121 82264
rect 57941 82180 57963 82236
rect 58019 82180 58043 82236
rect 58099 82180 58121 82236
rect 57941 82156 58121 82180
rect 57941 82100 57963 82156
rect 58019 82100 58043 82156
rect 58099 82100 58121 82156
rect 57941 82076 58121 82100
rect 57941 82020 57963 82076
rect 58019 82020 58043 82076
rect 58099 82020 58121 82076
rect 57941 81996 58121 82020
rect 57941 81940 57963 81996
rect 58019 81940 58043 81996
rect 58099 81940 58121 81996
rect 57941 81912 58121 81940
rect 59164 82236 59304 82264
rect 59164 82180 59206 82236
rect 59262 82180 59304 82236
rect 59164 82156 59304 82180
rect 59164 82100 59206 82156
rect 59262 82100 59304 82156
rect 59164 82076 59304 82100
rect 59164 82020 59206 82076
rect 59262 82020 59304 82076
rect 59164 81996 59304 82020
rect 59164 81940 59206 81996
rect 59262 81940 59304 81996
rect 59164 81912 59304 81940
rect 59334 82236 59450 82264
rect 59334 82180 59364 82236
rect 59420 82180 59450 82236
rect 59334 82156 59450 82180
rect 59334 82100 59364 82156
rect 59420 82100 59450 82156
rect 59334 82076 59450 82100
rect 59334 82020 59364 82076
rect 59420 82020 59450 82076
rect 59334 81996 59450 82020
rect 59334 81940 59364 81996
rect 59420 81940 59450 81996
rect 59334 81912 59450 81940
rect 59642 82236 59758 82264
rect 59642 82180 59672 82236
rect 59728 82180 59758 82236
rect 59642 82156 59758 82180
rect 59642 82100 59672 82156
rect 59728 82100 59758 82156
rect 59642 82076 59758 82100
rect 59642 82020 59672 82076
rect 59728 82020 59758 82076
rect 59642 81996 59758 82020
rect 59642 81940 59672 81996
rect 59728 81940 59758 81996
rect 59642 81912 59758 81940
rect 59788 82236 59904 82264
rect 59788 82180 59818 82236
rect 59874 82180 59904 82236
rect 59788 82156 59904 82180
rect 59788 82100 59818 82156
rect 59874 82100 59904 82156
rect 59788 82076 59904 82100
rect 59788 82020 59818 82076
rect 59874 82020 59904 82076
rect 59788 81996 59904 82020
rect 59788 81940 59818 81996
rect 59874 81940 59904 81996
rect 59788 81912 59904 81940
rect 59934 82236 60110 82264
rect 59934 82180 59954 82236
rect 60010 82180 60034 82236
rect 60090 82180 60110 82236
rect 59934 82156 60110 82180
rect 59934 82100 59954 82156
rect 60010 82100 60034 82156
rect 60090 82100 60110 82156
rect 59934 82076 60110 82100
rect 59934 82020 59954 82076
rect 60010 82020 60034 82076
rect 60090 82020 60110 82076
rect 59934 81996 60110 82020
rect 59934 81940 59954 81996
rect 60010 81940 60034 81996
rect 60090 81940 60110 81996
rect 59934 81912 60110 81940
rect 62307 82236 62481 82264
rect 62307 82180 62326 82236
rect 62382 82180 62406 82236
rect 62462 82180 62481 82236
rect 62307 82156 62481 82180
rect 62307 82100 62326 82156
rect 62382 82100 62406 82156
rect 62462 82100 62481 82156
rect 62307 82076 62481 82100
rect 62307 82020 62326 82076
rect 62382 82020 62406 82076
rect 62462 82020 62481 82076
rect 62307 81996 62481 82020
rect 62307 81940 62326 81996
rect 62382 81940 62406 81996
rect 62462 81940 62481 81996
rect 62307 81912 62481 81940
rect 64892 81802 64920 84186
rect 71836 83258 72188 84294
rect 71836 83206 71858 83258
rect 71910 83206 71922 83258
rect 71974 83206 71986 83258
rect 72038 83206 72050 83258
rect 72102 83206 72114 83258
rect 72166 83206 72188 83258
rect 65708 83156 65760 83162
rect 65708 83098 65760 83104
rect 64880 81796 64932 81802
rect 64880 81738 64932 81744
rect 64892 79898 64920 81738
rect 65524 80980 65576 80986
rect 65524 80922 65576 80928
rect 64880 79892 64932 79898
rect 64880 79834 64932 79840
rect 64892 77722 64920 79834
rect 64880 77716 64932 77722
rect 64880 77658 64932 77664
rect 64892 75206 64920 77658
rect 65340 76560 65392 76566
rect 65340 76502 65392 76508
rect 64880 75200 64932 75206
rect 64880 75142 64932 75148
rect 2020 74588 2124 74616
rect 2020 74532 2044 74588
rect 2100 74532 2124 74588
rect 2020 74508 2124 74532
rect 2020 74452 2044 74508
rect 2100 74452 2124 74508
rect 2020 74428 2124 74452
rect 2020 74372 2044 74428
rect 2100 74372 2124 74428
rect 2020 74348 2124 74372
rect 2020 74292 2044 74348
rect 2100 74292 2124 74348
rect 2020 74264 2124 74292
rect 5521 74588 5615 74616
rect 5521 74532 5540 74588
rect 5596 74532 5615 74588
rect 5521 74508 5615 74532
rect 5521 74452 5540 74508
rect 5596 74452 5615 74508
rect 5521 74428 5615 74452
rect 5521 74372 5540 74428
rect 5596 74372 5615 74428
rect 5521 74348 5615 74372
rect 5521 74292 5540 74348
rect 5596 74292 5615 74348
rect 5521 74264 5615 74292
rect 8411 74588 8505 74616
rect 8411 74532 8430 74588
rect 8486 74532 8505 74588
rect 8411 74508 8505 74532
rect 8411 74452 8430 74508
rect 8486 74452 8505 74508
rect 8411 74428 8505 74452
rect 8411 74372 8430 74428
rect 8486 74372 8505 74428
rect 8411 74348 8505 74372
rect 8411 74292 8430 74348
rect 8486 74292 8505 74348
rect 8411 74264 8505 74292
rect 11301 74588 11395 74616
rect 11301 74532 11320 74588
rect 11376 74532 11395 74588
rect 11301 74508 11395 74532
rect 11301 74452 11320 74508
rect 11376 74452 11395 74508
rect 11301 74428 11395 74452
rect 11301 74372 11320 74428
rect 11376 74372 11395 74428
rect 11301 74348 11395 74372
rect 11301 74292 11320 74348
rect 11376 74292 11395 74348
rect 11301 74264 11395 74292
rect 14191 74588 14285 74616
rect 14191 74532 14210 74588
rect 14266 74532 14285 74588
rect 14191 74508 14285 74532
rect 14191 74452 14210 74508
rect 14266 74452 14285 74508
rect 14191 74428 14285 74452
rect 14191 74372 14210 74428
rect 14266 74372 14285 74428
rect 14191 74348 14285 74372
rect 14191 74292 14210 74348
rect 14266 74292 14285 74348
rect 14191 74264 14285 74292
rect 17081 74588 17175 74616
rect 17081 74532 17100 74588
rect 17156 74532 17175 74588
rect 17081 74508 17175 74532
rect 17081 74452 17100 74508
rect 17156 74452 17175 74508
rect 17081 74428 17175 74452
rect 17081 74372 17100 74428
rect 17156 74372 17175 74428
rect 17081 74348 17175 74372
rect 17081 74292 17100 74348
rect 17156 74292 17175 74348
rect 17081 74264 17175 74292
rect 19971 74588 20065 74616
rect 19971 74532 19990 74588
rect 20046 74532 20065 74588
rect 19971 74508 20065 74532
rect 19971 74452 19990 74508
rect 20046 74452 20065 74508
rect 19971 74428 20065 74452
rect 19971 74372 19990 74428
rect 20046 74372 20065 74428
rect 19971 74348 20065 74372
rect 19971 74292 19990 74348
rect 20046 74292 20065 74348
rect 19971 74264 20065 74292
rect 22861 74588 22955 74616
rect 22861 74532 22880 74588
rect 22936 74532 22955 74588
rect 22861 74508 22955 74532
rect 22861 74452 22880 74508
rect 22936 74452 22955 74508
rect 22861 74428 22955 74452
rect 22861 74372 22880 74428
rect 22936 74372 22955 74428
rect 22861 74348 22955 74372
rect 22861 74292 22880 74348
rect 22936 74292 22955 74348
rect 22861 74264 22955 74292
rect 25751 74588 25845 74616
rect 25751 74532 25770 74588
rect 25826 74532 25845 74588
rect 25751 74508 25845 74532
rect 25751 74452 25770 74508
rect 25826 74452 25845 74508
rect 25751 74428 25845 74452
rect 25751 74372 25770 74428
rect 25826 74372 25845 74428
rect 25751 74348 25845 74372
rect 25751 74292 25770 74348
rect 25826 74292 25845 74348
rect 25751 74264 25845 74292
rect 28641 74588 28735 74616
rect 28641 74532 28660 74588
rect 28716 74532 28735 74588
rect 28641 74508 28735 74532
rect 28641 74452 28660 74508
rect 28716 74452 28735 74508
rect 28641 74428 28735 74452
rect 28641 74372 28660 74428
rect 28716 74372 28735 74428
rect 28641 74348 28735 74372
rect 28641 74292 28660 74348
rect 28716 74292 28735 74348
rect 28641 74264 28735 74292
rect 31531 74588 31625 74616
rect 31531 74532 31550 74588
rect 31606 74532 31625 74588
rect 31531 74508 31625 74532
rect 31531 74452 31550 74508
rect 31606 74452 31625 74508
rect 31531 74428 31625 74452
rect 31531 74372 31550 74428
rect 31606 74372 31625 74428
rect 31531 74348 31625 74372
rect 31531 74292 31550 74348
rect 31606 74292 31625 74348
rect 31531 74264 31625 74292
rect 34421 74588 34515 74616
rect 34421 74532 34440 74588
rect 34496 74532 34515 74588
rect 34421 74508 34515 74532
rect 34421 74452 34440 74508
rect 34496 74452 34515 74508
rect 34421 74428 34515 74452
rect 34421 74372 34440 74428
rect 34496 74372 34515 74428
rect 34421 74348 34515 74372
rect 34421 74292 34440 74348
rect 34496 74292 34515 74348
rect 34421 74264 34515 74292
rect 37311 74588 37405 74616
rect 37311 74532 37330 74588
rect 37386 74532 37405 74588
rect 37311 74508 37405 74532
rect 37311 74452 37330 74508
rect 37386 74452 37405 74508
rect 37311 74428 37405 74452
rect 37311 74372 37330 74428
rect 37386 74372 37405 74428
rect 37311 74348 37405 74372
rect 37311 74292 37330 74348
rect 37386 74292 37405 74348
rect 37311 74264 37405 74292
rect 40201 74588 40295 74616
rect 40201 74532 40220 74588
rect 40276 74532 40295 74588
rect 40201 74508 40295 74532
rect 40201 74452 40220 74508
rect 40276 74452 40295 74508
rect 40201 74428 40295 74452
rect 40201 74372 40220 74428
rect 40276 74372 40295 74428
rect 40201 74348 40295 74372
rect 40201 74292 40220 74348
rect 40276 74292 40295 74348
rect 40201 74264 40295 74292
rect 43091 74588 43185 74616
rect 43091 74532 43110 74588
rect 43166 74532 43185 74588
rect 43091 74508 43185 74532
rect 43091 74452 43110 74508
rect 43166 74452 43185 74508
rect 43091 74428 43185 74452
rect 43091 74372 43110 74428
rect 43166 74372 43185 74428
rect 43091 74348 43185 74372
rect 43091 74292 43110 74348
rect 43166 74292 43185 74348
rect 43091 74264 43185 74292
rect 45981 74588 46075 74616
rect 45981 74532 46000 74588
rect 46056 74532 46075 74588
rect 45981 74508 46075 74532
rect 45981 74452 46000 74508
rect 46056 74452 46075 74508
rect 45981 74428 46075 74452
rect 45981 74372 46000 74428
rect 46056 74372 46075 74428
rect 45981 74348 46075 74372
rect 45981 74292 46000 74348
rect 46056 74292 46075 74348
rect 45981 74264 46075 74292
rect 48989 74588 49083 74616
rect 48989 74532 49008 74588
rect 49064 74532 49083 74588
rect 48989 74508 49083 74532
rect 48989 74452 49008 74508
rect 49064 74452 49083 74508
rect 48989 74428 49083 74452
rect 48989 74372 49008 74428
rect 49064 74372 49083 74428
rect 48989 74348 49083 74372
rect 48989 74292 49008 74348
rect 49064 74292 49083 74348
rect 48989 74264 49083 74292
rect 52210 74588 52320 74616
rect 52210 74532 52237 74588
rect 52293 74532 52320 74588
rect 52210 74508 52320 74532
rect 52210 74452 52237 74508
rect 52293 74452 52320 74508
rect 52210 74428 52320 74452
rect 52210 74372 52237 74428
rect 52293 74372 52320 74428
rect 52210 74348 52320 74372
rect 52210 74292 52237 74348
rect 52293 74292 52320 74348
rect 52210 74264 52320 74292
rect 53602 74588 53730 74616
rect 53602 74532 53638 74588
rect 53694 74532 53730 74588
rect 53602 74508 53730 74532
rect 53602 74452 53638 74508
rect 53694 74452 53730 74508
rect 53602 74428 53730 74452
rect 53602 74372 53638 74428
rect 53694 74372 53730 74428
rect 53602 74348 53730 74372
rect 53602 74292 53638 74348
rect 53694 74292 53730 74348
rect 53602 74264 53730 74292
rect 53770 74588 53898 74616
rect 53770 74532 53806 74588
rect 53862 74532 53898 74588
rect 53770 74508 53898 74532
rect 53770 74452 53806 74508
rect 53862 74452 53898 74508
rect 53770 74428 53898 74452
rect 53770 74372 53806 74428
rect 53862 74372 53898 74428
rect 53770 74348 53898 74372
rect 53770 74292 53806 74348
rect 53862 74292 53898 74348
rect 53770 74264 53898 74292
rect 54514 74588 54642 74616
rect 54514 74532 54550 74588
rect 54606 74532 54642 74588
rect 54514 74508 54642 74532
rect 54514 74452 54550 74508
rect 54606 74452 54642 74508
rect 54514 74428 54642 74452
rect 54514 74372 54550 74428
rect 54606 74372 54642 74428
rect 54514 74348 54642 74372
rect 54514 74292 54550 74348
rect 54606 74292 54642 74348
rect 54514 74264 54642 74292
rect 54910 74588 55026 74616
rect 54910 74532 54940 74588
rect 54996 74532 55026 74588
rect 54910 74508 55026 74532
rect 54910 74452 54940 74508
rect 54996 74452 55026 74508
rect 54910 74428 55026 74452
rect 54910 74372 54940 74428
rect 54996 74372 55026 74428
rect 54910 74348 55026 74372
rect 54910 74292 54940 74348
rect 54996 74292 55026 74348
rect 54910 74264 55026 74292
rect 55620 74588 55748 74616
rect 55620 74532 55656 74588
rect 55712 74532 55748 74588
rect 55620 74508 55748 74532
rect 55620 74452 55656 74508
rect 55712 74452 55748 74508
rect 55620 74428 55748 74452
rect 55620 74372 55656 74428
rect 55712 74372 55748 74428
rect 55620 74348 55748 74372
rect 55620 74292 55656 74348
rect 55712 74292 55748 74348
rect 55620 74264 55748 74292
rect 56198 74588 56326 74616
rect 56198 74532 56234 74588
rect 56290 74532 56326 74588
rect 56198 74508 56326 74532
rect 56198 74452 56234 74508
rect 56290 74452 56326 74508
rect 56198 74428 56326 74452
rect 56198 74372 56234 74428
rect 56290 74372 56326 74428
rect 56198 74348 56326 74372
rect 56198 74292 56234 74348
rect 56290 74292 56326 74348
rect 56198 74264 56326 74292
rect 56649 74588 56765 74616
rect 56649 74532 56679 74588
rect 56735 74532 56765 74588
rect 56649 74508 56765 74532
rect 56649 74452 56679 74508
rect 56735 74452 56765 74508
rect 56649 74428 56765 74452
rect 56649 74372 56679 74428
rect 56735 74372 56765 74428
rect 56649 74348 56765 74372
rect 56649 74292 56679 74348
rect 56735 74292 56765 74348
rect 56649 74264 56765 74292
rect 56953 74588 57069 74616
rect 56953 74532 56983 74588
rect 57039 74532 57069 74588
rect 56953 74508 57069 74532
rect 56953 74452 56983 74508
rect 57039 74452 57069 74508
rect 56953 74428 57069 74452
rect 56953 74372 56983 74428
rect 57039 74372 57069 74428
rect 56953 74348 57069 74372
rect 56953 74292 56983 74348
rect 57039 74292 57069 74348
rect 56953 74264 57069 74292
rect 57795 74588 57911 74616
rect 57795 74532 57825 74588
rect 57881 74532 57911 74588
rect 57795 74508 57911 74532
rect 57795 74452 57825 74508
rect 57881 74452 57911 74508
rect 57795 74428 57911 74452
rect 57795 74372 57825 74428
rect 57881 74372 57911 74428
rect 57795 74348 57911 74372
rect 57795 74292 57825 74348
rect 57881 74292 57911 74348
rect 57795 74264 57911 74292
rect 58461 74588 58525 74616
rect 58461 74532 58465 74588
rect 58521 74532 58525 74588
rect 58461 74508 58525 74532
rect 58461 74452 58465 74508
rect 58521 74452 58525 74508
rect 58461 74428 58525 74452
rect 58461 74372 58465 74428
rect 58521 74372 58525 74428
rect 58461 74348 58525 74372
rect 58461 74292 58465 74348
rect 58521 74292 58525 74348
rect 58461 74264 58525 74292
rect 59018 74588 59134 74616
rect 59018 74532 59048 74588
rect 59104 74532 59134 74588
rect 59018 74508 59134 74532
rect 59018 74452 59048 74508
rect 59104 74452 59134 74508
rect 59018 74428 59134 74452
rect 59018 74372 59048 74428
rect 59104 74372 59134 74428
rect 59018 74348 59134 74372
rect 59018 74292 59048 74348
rect 59104 74292 59134 74348
rect 59018 74264 59134 74292
rect 60296 74588 60412 74616
rect 60296 74532 60326 74588
rect 60382 74532 60412 74588
rect 60296 74508 60412 74532
rect 60296 74452 60326 74508
rect 60382 74452 60412 74508
rect 60296 74428 60412 74452
rect 60296 74372 60326 74428
rect 60382 74372 60412 74428
rect 60296 74348 60412 74372
rect 60296 74292 60326 74348
rect 60382 74292 60412 74348
rect 60296 74264 60412 74292
rect 60454 74588 60570 74616
rect 60454 74532 60484 74588
rect 60540 74532 60570 74588
rect 60454 74508 60570 74532
rect 60454 74452 60484 74508
rect 60540 74452 60570 74508
rect 60454 74428 60570 74452
rect 60454 74372 60484 74428
rect 60540 74372 60570 74428
rect 60454 74348 60570 74372
rect 60454 74292 60484 74348
rect 60540 74292 60570 74348
rect 60454 74264 60570 74292
rect 62509 74588 62683 74616
rect 62509 74532 62528 74588
rect 62584 74532 62608 74588
rect 62664 74532 62683 74588
rect 62509 74508 62683 74532
rect 62509 74452 62528 74508
rect 62584 74452 62608 74508
rect 62664 74452 62683 74508
rect 62509 74428 62683 74452
rect 62509 74372 62528 74428
rect 62584 74372 62608 74428
rect 62664 74372 62683 74428
rect 62509 74348 62683 74372
rect 62509 74292 62528 74348
rect 62584 74292 62608 74348
rect 62664 74292 62683 74348
rect 62509 74264 62683 74292
rect 64892 73234 64920 75142
rect 64880 73228 64932 73234
rect 64880 73170 64932 73176
rect 2152 72236 2352 72264
rect 2152 72180 2184 72236
rect 2240 72180 2264 72236
rect 2320 72180 2352 72236
rect 2152 72156 2352 72180
rect 2152 72100 2184 72156
rect 2240 72100 2264 72156
rect 2320 72100 2352 72156
rect 2152 72076 2352 72100
rect 2152 72020 2184 72076
rect 2240 72020 2264 72076
rect 2320 72020 2352 72076
rect 2152 71996 2352 72020
rect 2152 71940 2184 71996
rect 2240 71940 2264 71996
rect 2320 71940 2352 71996
rect 2152 71912 2352 71940
rect 5374 72236 5468 72264
rect 5374 72180 5393 72236
rect 5449 72180 5468 72236
rect 5374 72156 5468 72180
rect 5374 72100 5393 72156
rect 5449 72100 5468 72156
rect 5374 72076 5468 72100
rect 5374 72020 5393 72076
rect 5449 72020 5468 72076
rect 5374 71996 5468 72020
rect 5374 71940 5393 71996
rect 5449 71940 5468 71996
rect 5374 71912 5468 71940
rect 8264 72236 8358 72264
rect 8264 72180 8283 72236
rect 8339 72180 8358 72236
rect 8264 72156 8358 72180
rect 8264 72100 8283 72156
rect 8339 72100 8358 72156
rect 8264 72076 8358 72100
rect 8264 72020 8283 72076
rect 8339 72020 8358 72076
rect 8264 71996 8358 72020
rect 8264 71940 8283 71996
rect 8339 71940 8358 71996
rect 8264 71912 8358 71940
rect 11154 72236 11248 72264
rect 11154 72180 11173 72236
rect 11229 72180 11248 72236
rect 11154 72156 11248 72180
rect 11154 72100 11173 72156
rect 11229 72100 11248 72156
rect 11154 72076 11248 72100
rect 11154 72020 11173 72076
rect 11229 72020 11248 72076
rect 11154 71996 11248 72020
rect 11154 71940 11173 71996
rect 11229 71940 11248 71996
rect 11154 71912 11248 71940
rect 14044 72236 14138 72264
rect 14044 72180 14063 72236
rect 14119 72180 14138 72236
rect 14044 72156 14138 72180
rect 14044 72100 14063 72156
rect 14119 72100 14138 72156
rect 14044 72076 14138 72100
rect 14044 72020 14063 72076
rect 14119 72020 14138 72076
rect 14044 71996 14138 72020
rect 14044 71940 14063 71996
rect 14119 71940 14138 71996
rect 14044 71912 14138 71940
rect 16934 72236 17028 72264
rect 16934 72180 16953 72236
rect 17009 72180 17028 72236
rect 16934 72156 17028 72180
rect 16934 72100 16953 72156
rect 17009 72100 17028 72156
rect 16934 72076 17028 72100
rect 16934 72020 16953 72076
rect 17009 72020 17028 72076
rect 16934 71996 17028 72020
rect 16934 71940 16953 71996
rect 17009 71940 17028 71996
rect 16934 71912 17028 71940
rect 19824 72236 19918 72264
rect 19824 72180 19843 72236
rect 19899 72180 19918 72236
rect 19824 72156 19918 72180
rect 19824 72100 19843 72156
rect 19899 72100 19918 72156
rect 19824 72076 19918 72100
rect 19824 72020 19843 72076
rect 19899 72020 19918 72076
rect 19824 71996 19918 72020
rect 19824 71940 19843 71996
rect 19899 71940 19918 71996
rect 19824 71912 19918 71940
rect 22714 72236 22808 72264
rect 22714 72180 22733 72236
rect 22789 72180 22808 72236
rect 22714 72156 22808 72180
rect 22714 72100 22733 72156
rect 22789 72100 22808 72156
rect 22714 72076 22808 72100
rect 22714 72020 22733 72076
rect 22789 72020 22808 72076
rect 22714 71996 22808 72020
rect 22714 71940 22733 71996
rect 22789 71940 22808 71996
rect 22714 71912 22808 71940
rect 25604 72236 25698 72264
rect 25604 72180 25623 72236
rect 25679 72180 25698 72236
rect 25604 72156 25698 72180
rect 25604 72100 25623 72156
rect 25679 72100 25698 72156
rect 25604 72076 25698 72100
rect 25604 72020 25623 72076
rect 25679 72020 25698 72076
rect 25604 71996 25698 72020
rect 25604 71940 25623 71996
rect 25679 71940 25698 71996
rect 25604 71912 25698 71940
rect 28494 72236 28588 72264
rect 28494 72180 28513 72236
rect 28569 72180 28588 72236
rect 28494 72156 28588 72180
rect 28494 72100 28513 72156
rect 28569 72100 28588 72156
rect 28494 72076 28588 72100
rect 28494 72020 28513 72076
rect 28569 72020 28588 72076
rect 28494 71996 28588 72020
rect 28494 71940 28513 71996
rect 28569 71940 28588 71996
rect 28494 71912 28588 71940
rect 31384 72236 31478 72264
rect 31384 72180 31403 72236
rect 31459 72180 31478 72236
rect 31384 72156 31478 72180
rect 31384 72100 31403 72156
rect 31459 72100 31478 72156
rect 31384 72076 31478 72100
rect 31384 72020 31403 72076
rect 31459 72020 31478 72076
rect 31384 71996 31478 72020
rect 31384 71940 31403 71996
rect 31459 71940 31478 71996
rect 31384 71912 31478 71940
rect 34274 72236 34368 72264
rect 34274 72180 34293 72236
rect 34349 72180 34368 72236
rect 34274 72156 34368 72180
rect 34274 72100 34293 72156
rect 34349 72100 34368 72156
rect 34274 72076 34368 72100
rect 34274 72020 34293 72076
rect 34349 72020 34368 72076
rect 34274 71996 34368 72020
rect 34274 71940 34293 71996
rect 34349 71940 34368 71996
rect 34274 71912 34368 71940
rect 37164 72236 37258 72264
rect 37164 72180 37183 72236
rect 37239 72180 37258 72236
rect 37164 72156 37258 72180
rect 37164 72100 37183 72156
rect 37239 72100 37258 72156
rect 37164 72076 37258 72100
rect 37164 72020 37183 72076
rect 37239 72020 37258 72076
rect 37164 71996 37258 72020
rect 37164 71940 37183 71996
rect 37239 71940 37258 71996
rect 37164 71912 37258 71940
rect 40054 72236 40148 72264
rect 40054 72180 40073 72236
rect 40129 72180 40148 72236
rect 40054 72156 40148 72180
rect 40054 72100 40073 72156
rect 40129 72100 40148 72156
rect 40054 72076 40148 72100
rect 40054 72020 40073 72076
rect 40129 72020 40148 72076
rect 40054 71996 40148 72020
rect 40054 71940 40073 71996
rect 40129 71940 40148 71996
rect 40054 71912 40148 71940
rect 42944 72236 43038 72264
rect 42944 72180 42963 72236
rect 43019 72180 43038 72236
rect 42944 72156 43038 72180
rect 42944 72100 42963 72156
rect 43019 72100 43038 72156
rect 42944 72076 43038 72100
rect 42944 72020 42963 72076
rect 43019 72020 43038 72076
rect 42944 71996 43038 72020
rect 42944 71940 42963 71996
rect 43019 71940 43038 71996
rect 42944 71912 43038 71940
rect 45834 72236 45928 72264
rect 45834 72180 45853 72236
rect 45909 72180 45928 72236
rect 45834 72156 45928 72180
rect 45834 72100 45853 72156
rect 45909 72100 45928 72156
rect 45834 72076 45928 72100
rect 45834 72020 45853 72076
rect 45909 72020 45928 72076
rect 45834 71996 45928 72020
rect 45834 71940 45853 71996
rect 45909 71940 45928 71996
rect 45834 71912 45928 71940
rect 48781 72236 48875 72264
rect 48781 72180 48800 72236
rect 48856 72180 48875 72236
rect 48781 72156 48875 72180
rect 48781 72100 48800 72156
rect 48856 72100 48875 72156
rect 48781 72076 48875 72100
rect 48781 72020 48800 72076
rect 48856 72020 48875 72076
rect 48781 71996 48875 72020
rect 48781 71940 48800 71996
rect 48856 71940 48875 71996
rect 48781 71912 48875 71940
rect 49630 72236 49830 72264
rect 49630 72180 49662 72236
rect 49718 72180 49742 72236
rect 49798 72180 49830 72236
rect 49630 72156 49830 72180
rect 49630 72100 49662 72156
rect 49718 72100 49742 72156
rect 49798 72100 49830 72156
rect 49630 72076 49830 72100
rect 49630 72020 49662 72076
rect 49718 72020 49742 72076
rect 49798 72020 49830 72076
rect 49630 71996 49830 72020
rect 49630 71940 49662 71996
rect 49718 71940 49742 71996
rect 49798 71940 49830 71996
rect 49630 71912 49830 71940
rect 52920 72236 53048 72264
rect 52920 72180 52956 72236
rect 53012 72180 53048 72236
rect 52920 72156 53048 72180
rect 52920 72100 52956 72156
rect 53012 72100 53048 72156
rect 52920 72076 53048 72100
rect 52920 72020 52956 72076
rect 53012 72020 53048 72076
rect 52920 71996 53048 72020
rect 52920 71940 52956 71996
rect 53012 71940 53048 71996
rect 52920 71912 53048 71940
rect 53078 72236 53206 72264
rect 53078 72180 53114 72236
rect 53170 72180 53206 72236
rect 53078 72156 53206 72180
rect 53078 72100 53114 72156
rect 53170 72100 53206 72156
rect 53078 72076 53206 72100
rect 53078 72020 53114 72076
rect 53170 72020 53206 72076
rect 53078 71996 53206 72020
rect 53078 71940 53114 71996
rect 53170 71940 53206 71996
rect 53078 71912 53206 71940
rect 53434 72236 53562 72264
rect 53434 72180 53470 72236
rect 53526 72180 53562 72236
rect 53434 72156 53562 72180
rect 53434 72100 53470 72156
rect 53526 72100 53562 72156
rect 53434 72076 53562 72100
rect 53434 72020 53470 72076
rect 53526 72020 53562 72076
rect 53434 71996 53562 72020
rect 53434 71940 53470 71996
rect 53526 71940 53562 71996
rect 53434 71912 53562 71940
rect 54752 72236 54880 72264
rect 54752 72180 54788 72236
rect 54844 72180 54880 72236
rect 54752 72156 54880 72180
rect 54752 72100 54788 72156
rect 54844 72100 54880 72156
rect 54752 72076 54880 72100
rect 54752 72020 54788 72076
rect 54844 72020 54880 72076
rect 54752 71996 54880 72020
rect 54752 71940 54788 71996
rect 54844 71940 54880 71996
rect 54752 71912 54880 71940
rect 55345 72236 55473 72264
rect 55345 72180 55381 72236
rect 55437 72180 55473 72236
rect 55345 72156 55473 72180
rect 55345 72100 55381 72156
rect 55437 72100 55473 72156
rect 55345 72076 55473 72100
rect 55345 72020 55381 72076
rect 55437 72020 55473 72076
rect 55345 71996 55473 72020
rect 55345 71940 55381 71996
rect 55437 71940 55473 71996
rect 55345 71912 55473 71940
rect 56491 72236 56619 72264
rect 56491 72180 56527 72236
rect 56583 72180 56619 72236
rect 56491 72156 56619 72180
rect 56491 72100 56527 72156
rect 56583 72100 56619 72156
rect 56491 72076 56619 72100
rect 56491 72020 56527 72076
rect 56583 72020 56619 72076
rect 56491 71996 56619 72020
rect 56491 71940 56527 71996
rect 56583 71940 56619 71996
rect 56491 71912 56619 71940
rect 57941 72236 58121 72264
rect 57941 72180 57963 72236
rect 58019 72180 58043 72236
rect 58099 72180 58121 72236
rect 57941 72156 58121 72180
rect 57941 72100 57963 72156
rect 58019 72100 58043 72156
rect 58099 72100 58121 72156
rect 57941 72076 58121 72100
rect 57941 72020 57963 72076
rect 58019 72020 58043 72076
rect 58099 72020 58121 72076
rect 57941 71996 58121 72020
rect 57941 71940 57963 71996
rect 58019 71940 58043 71996
rect 58099 71940 58121 71996
rect 57941 71912 58121 71940
rect 59164 72236 59304 72264
rect 59164 72180 59206 72236
rect 59262 72180 59304 72236
rect 59164 72156 59304 72180
rect 59164 72100 59206 72156
rect 59262 72100 59304 72156
rect 59164 72076 59304 72100
rect 59164 72020 59206 72076
rect 59262 72020 59304 72076
rect 59164 71996 59304 72020
rect 59164 71940 59206 71996
rect 59262 71940 59304 71996
rect 59164 71912 59304 71940
rect 59334 72236 59450 72264
rect 59334 72180 59364 72236
rect 59420 72180 59450 72236
rect 59334 72156 59450 72180
rect 59334 72100 59364 72156
rect 59420 72100 59450 72156
rect 59334 72076 59450 72100
rect 59334 72020 59364 72076
rect 59420 72020 59450 72076
rect 59334 71996 59450 72020
rect 59334 71940 59364 71996
rect 59420 71940 59450 71996
rect 59334 71912 59450 71940
rect 59642 72236 59758 72264
rect 59642 72180 59672 72236
rect 59728 72180 59758 72236
rect 59642 72156 59758 72180
rect 59642 72100 59672 72156
rect 59728 72100 59758 72156
rect 59642 72076 59758 72100
rect 59642 72020 59672 72076
rect 59728 72020 59758 72076
rect 59642 71996 59758 72020
rect 59642 71940 59672 71996
rect 59728 71940 59758 71996
rect 59642 71912 59758 71940
rect 59788 72236 59904 72264
rect 59788 72180 59818 72236
rect 59874 72180 59904 72236
rect 59788 72156 59904 72180
rect 59788 72100 59818 72156
rect 59874 72100 59904 72156
rect 59788 72076 59904 72100
rect 59788 72020 59818 72076
rect 59874 72020 59904 72076
rect 59788 71996 59904 72020
rect 59788 71940 59818 71996
rect 59874 71940 59904 71996
rect 59788 71912 59904 71940
rect 59934 72236 60110 72264
rect 59934 72180 59954 72236
rect 60010 72180 60034 72236
rect 60090 72180 60110 72236
rect 59934 72156 60110 72180
rect 59934 72100 59954 72156
rect 60010 72100 60034 72156
rect 60090 72100 60110 72156
rect 59934 72076 60110 72100
rect 59934 72020 59954 72076
rect 60010 72020 60034 72076
rect 60090 72020 60110 72076
rect 59934 71996 60110 72020
rect 59934 71940 59954 71996
rect 60010 71940 60034 71996
rect 60090 71940 60110 71996
rect 59934 71912 60110 71940
rect 62307 72236 62481 72264
rect 62307 72180 62326 72236
rect 62382 72180 62406 72236
rect 62462 72180 62481 72236
rect 62307 72156 62481 72180
rect 62307 72100 62326 72156
rect 62382 72100 62406 72156
rect 62462 72100 62481 72156
rect 62307 72076 62481 72100
rect 62307 72020 62326 72076
rect 62382 72020 62406 72076
rect 62462 72020 62481 72076
rect 62307 71996 62481 72020
rect 62307 71940 62326 71996
rect 62382 71940 62406 71996
rect 62462 71940 62481 71996
rect 62307 71912 62481 71940
rect 64604 71800 64656 71806
rect 64604 71742 64656 71748
rect 2020 64588 2124 64616
rect 2020 64532 2044 64588
rect 2100 64532 2124 64588
rect 2020 64508 2124 64532
rect 2020 64452 2044 64508
rect 2100 64452 2124 64508
rect 2020 64428 2124 64452
rect 2020 64372 2044 64428
rect 2100 64372 2124 64428
rect 2020 64348 2124 64372
rect 2020 64292 2044 64348
rect 2100 64292 2124 64348
rect 2020 64264 2124 64292
rect 5521 64588 5615 64616
rect 5521 64532 5540 64588
rect 5596 64532 5615 64588
rect 5521 64508 5615 64532
rect 5521 64452 5540 64508
rect 5596 64452 5615 64508
rect 5521 64428 5615 64452
rect 5521 64372 5540 64428
rect 5596 64372 5615 64428
rect 5521 64348 5615 64372
rect 5521 64292 5540 64348
rect 5596 64292 5615 64348
rect 5521 64264 5615 64292
rect 8411 64588 8505 64616
rect 8411 64532 8430 64588
rect 8486 64532 8505 64588
rect 8411 64508 8505 64532
rect 8411 64452 8430 64508
rect 8486 64452 8505 64508
rect 8411 64428 8505 64452
rect 8411 64372 8430 64428
rect 8486 64372 8505 64428
rect 8411 64348 8505 64372
rect 8411 64292 8430 64348
rect 8486 64292 8505 64348
rect 8411 64264 8505 64292
rect 11301 64588 11395 64616
rect 11301 64532 11320 64588
rect 11376 64532 11395 64588
rect 11301 64508 11395 64532
rect 11301 64452 11320 64508
rect 11376 64452 11395 64508
rect 11301 64428 11395 64452
rect 11301 64372 11320 64428
rect 11376 64372 11395 64428
rect 11301 64348 11395 64372
rect 11301 64292 11320 64348
rect 11376 64292 11395 64348
rect 11301 64264 11395 64292
rect 14191 64588 14285 64616
rect 14191 64532 14210 64588
rect 14266 64532 14285 64588
rect 14191 64508 14285 64532
rect 14191 64452 14210 64508
rect 14266 64452 14285 64508
rect 14191 64428 14285 64452
rect 14191 64372 14210 64428
rect 14266 64372 14285 64428
rect 14191 64348 14285 64372
rect 14191 64292 14210 64348
rect 14266 64292 14285 64348
rect 14191 64264 14285 64292
rect 17081 64588 17175 64616
rect 17081 64532 17100 64588
rect 17156 64532 17175 64588
rect 17081 64508 17175 64532
rect 17081 64452 17100 64508
rect 17156 64452 17175 64508
rect 17081 64428 17175 64452
rect 17081 64372 17100 64428
rect 17156 64372 17175 64428
rect 17081 64348 17175 64372
rect 17081 64292 17100 64348
rect 17156 64292 17175 64348
rect 17081 64264 17175 64292
rect 19971 64588 20065 64616
rect 19971 64532 19990 64588
rect 20046 64532 20065 64588
rect 19971 64508 20065 64532
rect 19971 64452 19990 64508
rect 20046 64452 20065 64508
rect 19971 64428 20065 64452
rect 19971 64372 19990 64428
rect 20046 64372 20065 64428
rect 19971 64348 20065 64372
rect 19971 64292 19990 64348
rect 20046 64292 20065 64348
rect 19971 64264 20065 64292
rect 22861 64588 22955 64616
rect 22861 64532 22880 64588
rect 22936 64532 22955 64588
rect 22861 64508 22955 64532
rect 22861 64452 22880 64508
rect 22936 64452 22955 64508
rect 22861 64428 22955 64452
rect 22861 64372 22880 64428
rect 22936 64372 22955 64428
rect 22861 64348 22955 64372
rect 22861 64292 22880 64348
rect 22936 64292 22955 64348
rect 22861 64264 22955 64292
rect 25751 64588 25845 64616
rect 25751 64532 25770 64588
rect 25826 64532 25845 64588
rect 25751 64508 25845 64532
rect 25751 64452 25770 64508
rect 25826 64452 25845 64508
rect 25751 64428 25845 64452
rect 25751 64372 25770 64428
rect 25826 64372 25845 64428
rect 25751 64348 25845 64372
rect 25751 64292 25770 64348
rect 25826 64292 25845 64348
rect 25751 64264 25845 64292
rect 28641 64588 28735 64616
rect 28641 64532 28660 64588
rect 28716 64532 28735 64588
rect 28641 64508 28735 64532
rect 28641 64452 28660 64508
rect 28716 64452 28735 64508
rect 28641 64428 28735 64452
rect 28641 64372 28660 64428
rect 28716 64372 28735 64428
rect 28641 64348 28735 64372
rect 28641 64292 28660 64348
rect 28716 64292 28735 64348
rect 28641 64264 28735 64292
rect 31531 64588 31625 64616
rect 31531 64532 31550 64588
rect 31606 64532 31625 64588
rect 31531 64508 31625 64532
rect 31531 64452 31550 64508
rect 31606 64452 31625 64508
rect 31531 64428 31625 64452
rect 31531 64372 31550 64428
rect 31606 64372 31625 64428
rect 31531 64348 31625 64372
rect 31531 64292 31550 64348
rect 31606 64292 31625 64348
rect 31531 64264 31625 64292
rect 34421 64588 34515 64616
rect 34421 64532 34440 64588
rect 34496 64532 34515 64588
rect 34421 64508 34515 64532
rect 34421 64452 34440 64508
rect 34496 64452 34515 64508
rect 34421 64428 34515 64452
rect 34421 64372 34440 64428
rect 34496 64372 34515 64428
rect 34421 64348 34515 64372
rect 34421 64292 34440 64348
rect 34496 64292 34515 64348
rect 34421 64264 34515 64292
rect 37311 64588 37405 64616
rect 37311 64532 37330 64588
rect 37386 64532 37405 64588
rect 37311 64508 37405 64532
rect 37311 64452 37330 64508
rect 37386 64452 37405 64508
rect 37311 64428 37405 64452
rect 37311 64372 37330 64428
rect 37386 64372 37405 64428
rect 37311 64348 37405 64372
rect 37311 64292 37330 64348
rect 37386 64292 37405 64348
rect 37311 64264 37405 64292
rect 40201 64588 40295 64616
rect 40201 64532 40220 64588
rect 40276 64532 40295 64588
rect 40201 64508 40295 64532
rect 40201 64452 40220 64508
rect 40276 64452 40295 64508
rect 40201 64428 40295 64452
rect 40201 64372 40220 64428
rect 40276 64372 40295 64428
rect 40201 64348 40295 64372
rect 40201 64292 40220 64348
rect 40276 64292 40295 64348
rect 40201 64264 40295 64292
rect 43091 64588 43185 64616
rect 43091 64532 43110 64588
rect 43166 64532 43185 64588
rect 43091 64508 43185 64532
rect 43091 64452 43110 64508
rect 43166 64452 43185 64508
rect 43091 64428 43185 64452
rect 43091 64372 43110 64428
rect 43166 64372 43185 64428
rect 43091 64348 43185 64372
rect 43091 64292 43110 64348
rect 43166 64292 43185 64348
rect 43091 64264 43185 64292
rect 45981 64588 46075 64616
rect 45981 64532 46000 64588
rect 46056 64532 46075 64588
rect 45981 64508 46075 64532
rect 45981 64452 46000 64508
rect 46056 64452 46075 64508
rect 45981 64428 46075 64452
rect 45981 64372 46000 64428
rect 46056 64372 46075 64428
rect 45981 64348 46075 64372
rect 45981 64292 46000 64348
rect 46056 64292 46075 64348
rect 45981 64264 46075 64292
rect 48989 64588 49083 64616
rect 48989 64532 49008 64588
rect 49064 64532 49083 64588
rect 48989 64508 49083 64532
rect 48989 64452 49008 64508
rect 49064 64452 49083 64508
rect 48989 64428 49083 64452
rect 48989 64372 49008 64428
rect 49064 64372 49083 64428
rect 48989 64348 49083 64372
rect 48989 64292 49008 64348
rect 49064 64292 49083 64348
rect 48989 64264 49083 64292
rect 52210 64588 52320 64616
rect 52210 64532 52237 64588
rect 52293 64532 52320 64588
rect 52210 64508 52320 64532
rect 52210 64452 52237 64508
rect 52293 64452 52320 64508
rect 52210 64428 52320 64452
rect 52210 64372 52237 64428
rect 52293 64372 52320 64428
rect 52210 64348 52320 64372
rect 52210 64292 52237 64348
rect 52293 64292 52320 64348
rect 52210 64264 52320 64292
rect 53602 64588 53730 64616
rect 53602 64532 53638 64588
rect 53694 64532 53730 64588
rect 53602 64508 53730 64532
rect 53602 64452 53638 64508
rect 53694 64452 53730 64508
rect 53602 64428 53730 64452
rect 53602 64372 53638 64428
rect 53694 64372 53730 64428
rect 53602 64348 53730 64372
rect 53602 64292 53638 64348
rect 53694 64292 53730 64348
rect 53602 64264 53730 64292
rect 53770 64588 53898 64616
rect 53770 64532 53806 64588
rect 53862 64532 53898 64588
rect 53770 64508 53898 64532
rect 53770 64452 53806 64508
rect 53862 64452 53898 64508
rect 53770 64428 53898 64452
rect 53770 64372 53806 64428
rect 53862 64372 53898 64428
rect 53770 64348 53898 64372
rect 53770 64292 53806 64348
rect 53862 64292 53898 64348
rect 53770 64264 53898 64292
rect 54514 64588 54642 64616
rect 54514 64532 54550 64588
rect 54606 64532 54642 64588
rect 54514 64508 54642 64532
rect 54514 64452 54550 64508
rect 54606 64452 54642 64508
rect 54514 64428 54642 64452
rect 54514 64372 54550 64428
rect 54606 64372 54642 64428
rect 54514 64348 54642 64372
rect 54514 64292 54550 64348
rect 54606 64292 54642 64348
rect 54514 64264 54642 64292
rect 54910 64588 55026 64616
rect 54910 64532 54940 64588
rect 54996 64532 55026 64588
rect 54910 64508 55026 64532
rect 54910 64452 54940 64508
rect 54996 64452 55026 64508
rect 54910 64428 55026 64452
rect 54910 64372 54940 64428
rect 54996 64372 55026 64428
rect 54910 64348 55026 64372
rect 54910 64292 54940 64348
rect 54996 64292 55026 64348
rect 54910 64264 55026 64292
rect 55620 64588 55748 64616
rect 55620 64532 55656 64588
rect 55712 64532 55748 64588
rect 55620 64508 55748 64532
rect 55620 64452 55656 64508
rect 55712 64452 55748 64508
rect 55620 64428 55748 64452
rect 55620 64372 55656 64428
rect 55712 64372 55748 64428
rect 55620 64348 55748 64372
rect 55620 64292 55656 64348
rect 55712 64292 55748 64348
rect 55620 64264 55748 64292
rect 56198 64588 56326 64616
rect 56198 64532 56234 64588
rect 56290 64532 56326 64588
rect 56198 64508 56326 64532
rect 56198 64452 56234 64508
rect 56290 64452 56326 64508
rect 56198 64428 56326 64452
rect 56198 64372 56234 64428
rect 56290 64372 56326 64428
rect 56198 64348 56326 64372
rect 56198 64292 56234 64348
rect 56290 64292 56326 64348
rect 56198 64264 56326 64292
rect 56649 64588 56765 64616
rect 56649 64532 56679 64588
rect 56735 64532 56765 64588
rect 56649 64508 56765 64532
rect 56649 64452 56679 64508
rect 56735 64452 56765 64508
rect 56649 64428 56765 64452
rect 56649 64372 56679 64428
rect 56735 64372 56765 64428
rect 56649 64348 56765 64372
rect 56649 64292 56679 64348
rect 56735 64292 56765 64348
rect 56649 64264 56765 64292
rect 56953 64588 57069 64616
rect 56953 64532 56983 64588
rect 57039 64532 57069 64588
rect 56953 64508 57069 64532
rect 56953 64452 56983 64508
rect 57039 64452 57069 64508
rect 56953 64428 57069 64452
rect 56953 64372 56983 64428
rect 57039 64372 57069 64428
rect 56953 64348 57069 64372
rect 56953 64292 56983 64348
rect 57039 64292 57069 64348
rect 56953 64264 57069 64292
rect 57795 64588 57911 64616
rect 57795 64532 57825 64588
rect 57881 64532 57911 64588
rect 57795 64508 57911 64532
rect 57795 64452 57825 64508
rect 57881 64452 57911 64508
rect 57795 64428 57911 64452
rect 57795 64372 57825 64428
rect 57881 64372 57911 64428
rect 57795 64348 57911 64372
rect 57795 64292 57825 64348
rect 57881 64292 57911 64348
rect 57795 64264 57911 64292
rect 58461 64588 58525 64616
rect 58461 64532 58465 64588
rect 58521 64532 58525 64588
rect 58461 64508 58525 64532
rect 58461 64452 58465 64508
rect 58521 64452 58525 64508
rect 58461 64428 58525 64452
rect 58461 64372 58465 64428
rect 58521 64372 58525 64428
rect 58461 64348 58525 64372
rect 58461 64292 58465 64348
rect 58521 64292 58525 64348
rect 58461 64264 58525 64292
rect 59018 64588 59134 64616
rect 59018 64532 59048 64588
rect 59104 64532 59134 64588
rect 59018 64508 59134 64532
rect 59018 64452 59048 64508
rect 59104 64452 59134 64508
rect 59018 64428 59134 64452
rect 59018 64372 59048 64428
rect 59104 64372 59134 64428
rect 59018 64348 59134 64372
rect 59018 64292 59048 64348
rect 59104 64292 59134 64348
rect 59018 64264 59134 64292
rect 60296 64588 60412 64616
rect 60296 64532 60326 64588
rect 60382 64532 60412 64588
rect 60296 64508 60412 64532
rect 60296 64452 60326 64508
rect 60382 64452 60412 64508
rect 60296 64428 60412 64452
rect 60296 64372 60326 64428
rect 60382 64372 60412 64428
rect 60296 64348 60412 64372
rect 60296 64292 60326 64348
rect 60382 64292 60412 64348
rect 60296 64264 60412 64292
rect 60454 64588 60570 64616
rect 60454 64532 60484 64588
rect 60540 64532 60570 64588
rect 60454 64508 60570 64532
rect 60454 64452 60484 64508
rect 60540 64452 60570 64508
rect 60454 64428 60570 64452
rect 60454 64372 60484 64428
rect 60540 64372 60570 64428
rect 60454 64348 60570 64372
rect 60454 64292 60484 64348
rect 60540 64292 60570 64348
rect 60454 64264 60570 64292
rect 62509 64588 62683 64616
rect 62509 64532 62528 64588
rect 62584 64532 62608 64588
rect 62664 64532 62683 64588
rect 62509 64508 62683 64532
rect 62509 64452 62528 64508
rect 62584 64452 62608 64508
rect 62664 64452 62683 64508
rect 62509 64428 62683 64452
rect 62509 64372 62528 64428
rect 62584 64372 62608 64428
rect 62664 64372 62683 64428
rect 62509 64348 62683 64372
rect 62509 64292 62528 64348
rect 62584 64292 62608 64348
rect 62664 64292 62683 64348
rect 62509 64264 62683 64292
rect 63592 63096 63644 63102
rect 63592 63038 63644 63044
rect 2152 62236 2352 62264
rect 2152 62180 2184 62236
rect 2240 62180 2264 62236
rect 2320 62180 2352 62236
rect 2152 62156 2352 62180
rect 2152 62100 2184 62156
rect 2240 62100 2264 62156
rect 2320 62100 2352 62156
rect 2152 62076 2352 62100
rect 2152 62020 2184 62076
rect 2240 62020 2264 62076
rect 2320 62020 2352 62076
rect 2152 61996 2352 62020
rect 2152 61940 2184 61996
rect 2240 61940 2264 61996
rect 2320 61940 2352 61996
rect 2152 61912 2352 61940
rect 5374 62236 5468 62264
rect 5374 62180 5393 62236
rect 5449 62180 5468 62236
rect 5374 62156 5468 62180
rect 5374 62100 5393 62156
rect 5449 62100 5468 62156
rect 5374 62076 5468 62100
rect 5374 62020 5393 62076
rect 5449 62020 5468 62076
rect 5374 61996 5468 62020
rect 5374 61940 5393 61996
rect 5449 61940 5468 61996
rect 5374 61912 5468 61940
rect 8264 62236 8358 62264
rect 8264 62180 8283 62236
rect 8339 62180 8358 62236
rect 8264 62156 8358 62180
rect 8264 62100 8283 62156
rect 8339 62100 8358 62156
rect 8264 62076 8358 62100
rect 8264 62020 8283 62076
rect 8339 62020 8358 62076
rect 8264 61996 8358 62020
rect 8264 61940 8283 61996
rect 8339 61940 8358 61996
rect 8264 61912 8358 61940
rect 11154 62236 11248 62264
rect 11154 62180 11173 62236
rect 11229 62180 11248 62236
rect 11154 62156 11248 62180
rect 11154 62100 11173 62156
rect 11229 62100 11248 62156
rect 11154 62076 11248 62100
rect 11154 62020 11173 62076
rect 11229 62020 11248 62076
rect 11154 61996 11248 62020
rect 11154 61940 11173 61996
rect 11229 61940 11248 61996
rect 11154 61912 11248 61940
rect 14044 62236 14138 62264
rect 14044 62180 14063 62236
rect 14119 62180 14138 62236
rect 14044 62156 14138 62180
rect 14044 62100 14063 62156
rect 14119 62100 14138 62156
rect 14044 62076 14138 62100
rect 14044 62020 14063 62076
rect 14119 62020 14138 62076
rect 14044 61996 14138 62020
rect 14044 61940 14063 61996
rect 14119 61940 14138 61996
rect 14044 61912 14138 61940
rect 16934 62236 17028 62264
rect 16934 62180 16953 62236
rect 17009 62180 17028 62236
rect 16934 62156 17028 62180
rect 16934 62100 16953 62156
rect 17009 62100 17028 62156
rect 16934 62076 17028 62100
rect 16934 62020 16953 62076
rect 17009 62020 17028 62076
rect 16934 61996 17028 62020
rect 16934 61940 16953 61996
rect 17009 61940 17028 61996
rect 16934 61912 17028 61940
rect 19824 62236 19918 62264
rect 19824 62180 19843 62236
rect 19899 62180 19918 62236
rect 19824 62156 19918 62180
rect 19824 62100 19843 62156
rect 19899 62100 19918 62156
rect 19824 62076 19918 62100
rect 19824 62020 19843 62076
rect 19899 62020 19918 62076
rect 19824 61996 19918 62020
rect 19824 61940 19843 61996
rect 19899 61940 19918 61996
rect 19824 61912 19918 61940
rect 22714 62236 22808 62264
rect 22714 62180 22733 62236
rect 22789 62180 22808 62236
rect 22714 62156 22808 62180
rect 22714 62100 22733 62156
rect 22789 62100 22808 62156
rect 22714 62076 22808 62100
rect 22714 62020 22733 62076
rect 22789 62020 22808 62076
rect 22714 61996 22808 62020
rect 22714 61940 22733 61996
rect 22789 61940 22808 61996
rect 22714 61912 22808 61940
rect 25604 62236 25698 62264
rect 25604 62180 25623 62236
rect 25679 62180 25698 62236
rect 25604 62156 25698 62180
rect 25604 62100 25623 62156
rect 25679 62100 25698 62156
rect 25604 62076 25698 62100
rect 25604 62020 25623 62076
rect 25679 62020 25698 62076
rect 25604 61996 25698 62020
rect 25604 61940 25623 61996
rect 25679 61940 25698 61996
rect 25604 61912 25698 61940
rect 28494 62236 28588 62264
rect 28494 62180 28513 62236
rect 28569 62180 28588 62236
rect 28494 62156 28588 62180
rect 28494 62100 28513 62156
rect 28569 62100 28588 62156
rect 28494 62076 28588 62100
rect 28494 62020 28513 62076
rect 28569 62020 28588 62076
rect 28494 61996 28588 62020
rect 28494 61940 28513 61996
rect 28569 61940 28588 61996
rect 28494 61912 28588 61940
rect 31384 62236 31478 62264
rect 31384 62180 31403 62236
rect 31459 62180 31478 62236
rect 31384 62156 31478 62180
rect 31384 62100 31403 62156
rect 31459 62100 31478 62156
rect 31384 62076 31478 62100
rect 31384 62020 31403 62076
rect 31459 62020 31478 62076
rect 31384 61996 31478 62020
rect 31384 61940 31403 61996
rect 31459 61940 31478 61996
rect 31384 61912 31478 61940
rect 34274 62236 34368 62264
rect 34274 62180 34293 62236
rect 34349 62180 34368 62236
rect 34274 62156 34368 62180
rect 34274 62100 34293 62156
rect 34349 62100 34368 62156
rect 34274 62076 34368 62100
rect 34274 62020 34293 62076
rect 34349 62020 34368 62076
rect 34274 61996 34368 62020
rect 34274 61940 34293 61996
rect 34349 61940 34368 61996
rect 34274 61912 34368 61940
rect 37164 62236 37258 62264
rect 37164 62180 37183 62236
rect 37239 62180 37258 62236
rect 37164 62156 37258 62180
rect 37164 62100 37183 62156
rect 37239 62100 37258 62156
rect 37164 62076 37258 62100
rect 37164 62020 37183 62076
rect 37239 62020 37258 62076
rect 37164 61996 37258 62020
rect 37164 61940 37183 61996
rect 37239 61940 37258 61996
rect 37164 61912 37258 61940
rect 40054 62236 40148 62264
rect 40054 62180 40073 62236
rect 40129 62180 40148 62236
rect 40054 62156 40148 62180
rect 40054 62100 40073 62156
rect 40129 62100 40148 62156
rect 40054 62076 40148 62100
rect 40054 62020 40073 62076
rect 40129 62020 40148 62076
rect 40054 61996 40148 62020
rect 40054 61940 40073 61996
rect 40129 61940 40148 61996
rect 40054 61912 40148 61940
rect 42944 62236 43038 62264
rect 42944 62180 42963 62236
rect 43019 62180 43038 62236
rect 42944 62156 43038 62180
rect 42944 62100 42963 62156
rect 43019 62100 43038 62156
rect 42944 62076 43038 62100
rect 42944 62020 42963 62076
rect 43019 62020 43038 62076
rect 42944 61996 43038 62020
rect 42944 61940 42963 61996
rect 43019 61940 43038 61996
rect 42944 61912 43038 61940
rect 45834 62236 45928 62264
rect 45834 62180 45853 62236
rect 45909 62180 45928 62236
rect 45834 62156 45928 62180
rect 45834 62100 45853 62156
rect 45909 62100 45928 62156
rect 45834 62076 45928 62100
rect 45834 62020 45853 62076
rect 45909 62020 45928 62076
rect 45834 61996 45928 62020
rect 45834 61940 45853 61996
rect 45909 61940 45928 61996
rect 45834 61912 45928 61940
rect 48781 62236 48875 62264
rect 48781 62180 48800 62236
rect 48856 62180 48875 62236
rect 48781 62156 48875 62180
rect 48781 62100 48800 62156
rect 48856 62100 48875 62156
rect 48781 62076 48875 62100
rect 48781 62020 48800 62076
rect 48856 62020 48875 62076
rect 48781 61996 48875 62020
rect 48781 61940 48800 61996
rect 48856 61940 48875 61996
rect 48781 61912 48875 61940
rect 49630 62236 49830 62264
rect 49630 62180 49662 62236
rect 49718 62180 49742 62236
rect 49798 62180 49830 62236
rect 49630 62156 49830 62180
rect 49630 62100 49662 62156
rect 49718 62100 49742 62156
rect 49798 62100 49830 62156
rect 49630 62076 49830 62100
rect 49630 62020 49662 62076
rect 49718 62020 49742 62076
rect 49798 62020 49830 62076
rect 49630 61996 49830 62020
rect 49630 61940 49662 61996
rect 49718 61940 49742 61996
rect 49798 61940 49830 61996
rect 49630 61912 49830 61940
rect 52920 62236 53048 62264
rect 52920 62180 52956 62236
rect 53012 62180 53048 62236
rect 52920 62156 53048 62180
rect 52920 62100 52956 62156
rect 53012 62100 53048 62156
rect 52920 62076 53048 62100
rect 52920 62020 52956 62076
rect 53012 62020 53048 62076
rect 52920 61996 53048 62020
rect 52920 61940 52956 61996
rect 53012 61940 53048 61996
rect 52920 61912 53048 61940
rect 53078 62236 53206 62264
rect 53078 62180 53114 62236
rect 53170 62180 53206 62236
rect 53078 62156 53206 62180
rect 53078 62100 53114 62156
rect 53170 62100 53206 62156
rect 53078 62076 53206 62100
rect 53078 62020 53114 62076
rect 53170 62020 53206 62076
rect 53078 61996 53206 62020
rect 53078 61940 53114 61996
rect 53170 61940 53206 61996
rect 53078 61912 53206 61940
rect 53434 62236 53562 62264
rect 53434 62180 53470 62236
rect 53526 62180 53562 62236
rect 53434 62156 53562 62180
rect 53434 62100 53470 62156
rect 53526 62100 53562 62156
rect 53434 62076 53562 62100
rect 53434 62020 53470 62076
rect 53526 62020 53562 62076
rect 53434 61996 53562 62020
rect 53434 61940 53470 61996
rect 53526 61940 53562 61996
rect 53434 61912 53562 61940
rect 54752 62236 54880 62264
rect 54752 62180 54788 62236
rect 54844 62180 54880 62236
rect 54752 62156 54880 62180
rect 54752 62100 54788 62156
rect 54844 62100 54880 62156
rect 54752 62076 54880 62100
rect 54752 62020 54788 62076
rect 54844 62020 54880 62076
rect 54752 61996 54880 62020
rect 54752 61940 54788 61996
rect 54844 61940 54880 61996
rect 54752 61912 54880 61940
rect 55345 62236 55473 62264
rect 55345 62180 55381 62236
rect 55437 62180 55473 62236
rect 55345 62156 55473 62180
rect 55345 62100 55381 62156
rect 55437 62100 55473 62156
rect 55345 62076 55473 62100
rect 55345 62020 55381 62076
rect 55437 62020 55473 62076
rect 55345 61996 55473 62020
rect 55345 61940 55381 61996
rect 55437 61940 55473 61996
rect 55345 61912 55473 61940
rect 56491 62236 56619 62264
rect 56491 62180 56527 62236
rect 56583 62180 56619 62236
rect 56491 62156 56619 62180
rect 56491 62100 56527 62156
rect 56583 62100 56619 62156
rect 56491 62076 56619 62100
rect 56491 62020 56527 62076
rect 56583 62020 56619 62076
rect 56491 61996 56619 62020
rect 56491 61940 56527 61996
rect 56583 61940 56619 61996
rect 56491 61912 56619 61940
rect 57941 62236 58121 62264
rect 57941 62180 57963 62236
rect 58019 62180 58043 62236
rect 58099 62180 58121 62236
rect 57941 62156 58121 62180
rect 57941 62100 57963 62156
rect 58019 62100 58043 62156
rect 58099 62100 58121 62156
rect 57941 62076 58121 62100
rect 57941 62020 57963 62076
rect 58019 62020 58043 62076
rect 58099 62020 58121 62076
rect 57941 61996 58121 62020
rect 57941 61940 57963 61996
rect 58019 61940 58043 61996
rect 58099 61940 58121 61996
rect 57941 61912 58121 61940
rect 59164 62236 59304 62264
rect 59164 62180 59206 62236
rect 59262 62180 59304 62236
rect 59164 62156 59304 62180
rect 59164 62100 59206 62156
rect 59262 62100 59304 62156
rect 59164 62076 59304 62100
rect 59164 62020 59206 62076
rect 59262 62020 59304 62076
rect 59164 61996 59304 62020
rect 59164 61940 59206 61996
rect 59262 61940 59304 61996
rect 59164 61912 59304 61940
rect 59334 62236 59450 62264
rect 59334 62180 59364 62236
rect 59420 62180 59450 62236
rect 59334 62156 59450 62180
rect 59334 62100 59364 62156
rect 59420 62100 59450 62156
rect 59334 62076 59450 62100
rect 59334 62020 59364 62076
rect 59420 62020 59450 62076
rect 59334 61996 59450 62020
rect 59334 61940 59364 61996
rect 59420 61940 59450 61996
rect 59334 61912 59450 61940
rect 59642 62236 59758 62264
rect 59642 62180 59672 62236
rect 59728 62180 59758 62236
rect 59642 62156 59758 62180
rect 59642 62100 59672 62156
rect 59728 62100 59758 62156
rect 59642 62076 59758 62100
rect 59642 62020 59672 62076
rect 59728 62020 59758 62076
rect 59642 61996 59758 62020
rect 59642 61940 59672 61996
rect 59728 61940 59758 61996
rect 59642 61912 59758 61940
rect 59788 62236 59904 62264
rect 59788 62180 59818 62236
rect 59874 62180 59904 62236
rect 59788 62156 59904 62180
rect 59788 62100 59818 62156
rect 59874 62100 59904 62156
rect 59788 62076 59904 62100
rect 59788 62020 59818 62076
rect 59874 62020 59904 62076
rect 59788 61996 59904 62020
rect 59788 61940 59818 61996
rect 59874 61940 59904 61996
rect 59788 61912 59904 61940
rect 59934 62236 60110 62264
rect 59934 62180 59954 62236
rect 60010 62180 60034 62236
rect 60090 62180 60110 62236
rect 59934 62156 60110 62180
rect 59934 62100 59954 62156
rect 60010 62100 60034 62156
rect 60090 62100 60110 62156
rect 59934 62076 60110 62100
rect 59934 62020 59954 62076
rect 60010 62020 60034 62076
rect 60090 62020 60110 62076
rect 59934 61996 60110 62020
rect 59934 61940 59954 61996
rect 60010 61940 60034 61996
rect 60090 61940 60110 61996
rect 59934 61912 60110 61940
rect 62307 62236 62481 62264
rect 62307 62180 62326 62236
rect 62382 62180 62406 62236
rect 62462 62180 62481 62236
rect 62307 62156 62481 62180
rect 62307 62100 62326 62156
rect 62382 62100 62406 62156
rect 62462 62100 62481 62156
rect 62307 62076 62481 62100
rect 62307 62020 62326 62076
rect 62382 62020 62406 62076
rect 62462 62020 62481 62076
rect 62307 61996 62481 62020
rect 62307 61940 62326 61996
rect 62382 61940 62406 61996
rect 62462 61940 62481 61996
rect 62307 61912 62481 61940
rect 63500 61230 63552 61236
rect 63500 61172 63552 61178
rect 2020 54588 2124 54616
rect 2020 54532 2044 54588
rect 2100 54532 2124 54588
rect 2020 54508 2124 54532
rect 2020 54452 2044 54508
rect 2100 54452 2124 54508
rect 2020 54428 2124 54452
rect 2020 54372 2044 54428
rect 2100 54372 2124 54428
rect 2020 54348 2124 54372
rect 2020 54292 2044 54348
rect 2100 54292 2124 54348
rect 2020 54264 2124 54292
rect 5521 54588 5615 54616
rect 5521 54532 5540 54588
rect 5596 54532 5615 54588
rect 5521 54508 5615 54532
rect 5521 54452 5540 54508
rect 5596 54452 5615 54508
rect 5521 54428 5615 54452
rect 5521 54372 5540 54428
rect 5596 54372 5615 54428
rect 5521 54348 5615 54372
rect 5521 54292 5540 54348
rect 5596 54292 5615 54348
rect 5521 54264 5615 54292
rect 8411 54588 8505 54616
rect 8411 54532 8430 54588
rect 8486 54532 8505 54588
rect 8411 54508 8505 54532
rect 8411 54452 8430 54508
rect 8486 54452 8505 54508
rect 8411 54428 8505 54452
rect 8411 54372 8430 54428
rect 8486 54372 8505 54428
rect 8411 54348 8505 54372
rect 8411 54292 8430 54348
rect 8486 54292 8505 54348
rect 8411 54264 8505 54292
rect 11301 54588 11395 54616
rect 11301 54532 11320 54588
rect 11376 54532 11395 54588
rect 11301 54508 11395 54532
rect 11301 54452 11320 54508
rect 11376 54452 11395 54508
rect 11301 54428 11395 54452
rect 11301 54372 11320 54428
rect 11376 54372 11395 54428
rect 11301 54348 11395 54372
rect 11301 54292 11320 54348
rect 11376 54292 11395 54348
rect 11301 54264 11395 54292
rect 14191 54588 14285 54616
rect 14191 54532 14210 54588
rect 14266 54532 14285 54588
rect 14191 54508 14285 54532
rect 14191 54452 14210 54508
rect 14266 54452 14285 54508
rect 14191 54428 14285 54452
rect 14191 54372 14210 54428
rect 14266 54372 14285 54428
rect 14191 54348 14285 54372
rect 14191 54292 14210 54348
rect 14266 54292 14285 54348
rect 14191 54264 14285 54292
rect 17081 54588 17175 54616
rect 17081 54532 17100 54588
rect 17156 54532 17175 54588
rect 17081 54508 17175 54532
rect 17081 54452 17100 54508
rect 17156 54452 17175 54508
rect 17081 54428 17175 54452
rect 17081 54372 17100 54428
rect 17156 54372 17175 54428
rect 17081 54348 17175 54372
rect 17081 54292 17100 54348
rect 17156 54292 17175 54348
rect 17081 54264 17175 54292
rect 19971 54588 20065 54616
rect 19971 54532 19990 54588
rect 20046 54532 20065 54588
rect 19971 54508 20065 54532
rect 19971 54452 19990 54508
rect 20046 54452 20065 54508
rect 19971 54428 20065 54452
rect 19971 54372 19990 54428
rect 20046 54372 20065 54428
rect 19971 54348 20065 54372
rect 19971 54292 19990 54348
rect 20046 54292 20065 54348
rect 19971 54264 20065 54292
rect 22861 54588 22955 54616
rect 22861 54532 22880 54588
rect 22936 54532 22955 54588
rect 22861 54508 22955 54532
rect 22861 54452 22880 54508
rect 22936 54452 22955 54508
rect 22861 54428 22955 54452
rect 22861 54372 22880 54428
rect 22936 54372 22955 54428
rect 22861 54348 22955 54372
rect 22861 54292 22880 54348
rect 22936 54292 22955 54348
rect 22861 54264 22955 54292
rect 25751 54588 25845 54616
rect 25751 54532 25770 54588
rect 25826 54532 25845 54588
rect 25751 54508 25845 54532
rect 25751 54452 25770 54508
rect 25826 54452 25845 54508
rect 25751 54428 25845 54452
rect 25751 54372 25770 54428
rect 25826 54372 25845 54428
rect 25751 54348 25845 54372
rect 25751 54292 25770 54348
rect 25826 54292 25845 54348
rect 25751 54264 25845 54292
rect 28641 54588 28735 54616
rect 28641 54532 28660 54588
rect 28716 54532 28735 54588
rect 28641 54508 28735 54532
rect 28641 54452 28660 54508
rect 28716 54452 28735 54508
rect 28641 54428 28735 54452
rect 28641 54372 28660 54428
rect 28716 54372 28735 54428
rect 28641 54348 28735 54372
rect 28641 54292 28660 54348
rect 28716 54292 28735 54348
rect 28641 54264 28735 54292
rect 31531 54588 31625 54616
rect 31531 54532 31550 54588
rect 31606 54532 31625 54588
rect 31531 54508 31625 54532
rect 31531 54452 31550 54508
rect 31606 54452 31625 54508
rect 31531 54428 31625 54452
rect 31531 54372 31550 54428
rect 31606 54372 31625 54428
rect 31531 54348 31625 54372
rect 31531 54292 31550 54348
rect 31606 54292 31625 54348
rect 31531 54264 31625 54292
rect 34421 54588 34515 54616
rect 34421 54532 34440 54588
rect 34496 54532 34515 54588
rect 34421 54508 34515 54532
rect 34421 54452 34440 54508
rect 34496 54452 34515 54508
rect 34421 54428 34515 54452
rect 34421 54372 34440 54428
rect 34496 54372 34515 54428
rect 34421 54348 34515 54372
rect 34421 54292 34440 54348
rect 34496 54292 34515 54348
rect 34421 54264 34515 54292
rect 37311 54588 37405 54616
rect 37311 54532 37330 54588
rect 37386 54532 37405 54588
rect 37311 54508 37405 54532
rect 37311 54452 37330 54508
rect 37386 54452 37405 54508
rect 37311 54428 37405 54452
rect 37311 54372 37330 54428
rect 37386 54372 37405 54428
rect 37311 54348 37405 54372
rect 37311 54292 37330 54348
rect 37386 54292 37405 54348
rect 37311 54264 37405 54292
rect 40201 54588 40295 54616
rect 40201 54532 40220 54588
rect 40276 54532 40295 54588
rect 40201 54508 40295 54532
rect 40201 54452 40220 54508
rect 40276 54452 40295 54508
rect 40201 54428 40295 54452
rect 40201 54372 40220 54428
rect 40276 54372 40295 54428
rect 40201 54348 40295 54372
rect 40201 54292 40220 54348
rect 40276 54292 40295 54348
rect 40201 54264 40295 54292
rect 43091 54588 43185 54616
rect 43091 54532 43110 54588
rect 43166 54532 43185 54588
rect 43091 54508 43185 54532
rect 43091 54452 43110 54508
rect 43166 54452 43185 54508
rect 43091 54428 43185 54452
rect 43091 54372 43110 54428
rect 43166 54372 43185 54428
rect 43091 54348 43185 54372
rect 43091 54292 43110 54348
rect 43166 54292 43185 54348
rect 43091 54264 43185 54292
rect 45981 54588 46075 54616
rect 45981 54532 46000 54588
rect 46056 54532 46075 54588
rect 45981 54508 46075 54532
rect 45981 54452 46000 54508
rect 46056 54452 46075 54508
rect 45981 54428 46075 54452
rect 45981 54372 46000 54428
rect 46056 54372 46075 54428
rect 45981 54348 46075 54372
rect 45981 54292 46000 54348
rect 46056 54292 46075 54348
rect 45981 54264 46075 54292
rect 48989 54588 49083 54616
rect 48989 54532 49008 54588
rect 49064 54532 49083 54588
rect 48989 54508 49083 54532
rect 48989 54452 49008 54508
rect 49064 54452 49083 54508
rect 48989 54428 49083 54452
rect 48989 54372 49008 54428
rect 49064 54372 49083 54428
rect 48989 54348 49083 54372
rect 48989 54292 49008 54348
rect 49064 54292 49083 54348
rect 48989 54264 49083 54292
rect 52210 54588 52320 54616
rect 52210 54532 52237 54588
rect 52293 54532 52320 54588
rect 52210 54508 52320 54532
rect 52210 54452 52237 54508
rect 52293 54452 52320 54508
rect 52210 54428 52320 54452
rect 52210 54372 52237 54428
rect 52293 54372 52320 54428
rect 52210 54348 52320 54372
rect 52210 54292 52237 54348
rect 52293 54292 52320 54348
rect 52210 54264 52320 54292
rect 53602 54588 53730 54616
rect 53602 54532 53638 54588
rect 53694 54532 53730 54588
rect 53602 54508 53730 54532
rect 53602 54452 53638 54508
rect 53694 54452 53730 54508
rect 53602 54428 53730 54452
rect 53602 54372 53638 54428
rect 53694 54372 53730 54428
rect 53602 54348 53730 54372
rect 53602 54292 53638 54348
rect 53694 54292 53730 54348
rect 53602 54264 53730 54292
rect 53770 54588 53898 54616
rect 53770 54532 53806 54588
rect 53862 54532 53898 54588
rect 53770 54508 53898 54532
rect 53770 54452 53806 54508
rect 53862 54452 53898 54508
rect 53770 54428 53898 54452
rect 53770 54372 53806 54428
rect 53862 54372 53898 54428
rect 53770 54348 53898 54372
rect 53770 54292 53806 54348
rect 53862 54292 53898 54348
rect 53770 54264 53898 54292
rect 54514 54588 54642 54616
rect 54514 54532 54550 54588
rect 54606 54532 54642 54588
rect 54514 54508 54642 54532
rect 54514 54452 54550 54508
rect 54606 54452 54642 54508
rect 54514 54428 54642 54452
rect 54514 54372 54550 54428
rect 54606 54372 54642 54428
rect 54514 54348 54642 54372
rect 54514 54292 54550 54348
rect 54606 54292 54642 54348
rect 54514 54264 54642 54292
rect 54910 54588 55026 54616
rect 54910 54532 54940 54588
rect 54996 54532 55026 54588
rect 54910 54508 55026 54532
rect 54910 54452 54940 54508
rect 54996 54452 55026 54508
rect 54910 54428 55026 54452
rect 54910 54372 54940 54428
rect 54996 54372 55026 54428
rect 54910 54348 55026 54372
rect 54910 54292 54940 54348
rect 54996 54292 55026 54348
rect 54910 54264 55026 54292
rect 55620 54588 55748 54616
rect 55620 54532 55656 54588
rect 55712 54532 55748 54588
rect 55620 54508 55748 54532
rect 55620 54452 55656 54508
rect 55712 54452 55748 54508
rect 55620 54428 55748 54452
rect 55620 54372 55656 54428
rect 55712 54372 55748 54428
rect 55620 54348 55748 54372
rect 55620 54292 55656 54348
rect 55712 54292 55748 54348
rect 55620 54264 55748 54292
rect 56198 54588 56326 54616
rect 56198 54532 56234 54588
rect 56290 54532 56326 54588
rect 56198 54508 56326 54532
rect 56198 54452 56234 54508
rect 56290 54452 56326 54508
rect 56198 54428 56326 54452
rect 56198 54372 56234 54428
rect 56290 54372 56326 54428
rect 56198 54348 56326 54372
rect 56198 54292 56234 54348
rect 56290 54292 56326 54348
rect 56198 54264 56326 54292
rect 56649 54588 56765 54616
rect 56649 54532 56679 54588
rect 56735 54532 56765 54588
rect 56649 54508 56765 54532
rect 56649 54452 56679 54508
rect 56735 54452 56765 54508
rect 56649 54428 56765 54452
rect 56649 54372 56679 54428
rect 56735 54372 56765 54428
rect 56649 54348 56765 54372
rect 56649 54292 56679 54348
rect 56735 54292 56765 54348
rect 56649 54264 56765 54292
rect 56953 54588 57069 54616
rect 56953 54532 56983 54588
rect 57039 54532 57069 54588
rect 56953 54508 57069 54532
rect 56953 54452 56983 54508
rect 57039 54452 57069 54508
rect 56953 54428 57069 54452
rect 56953 54372 56983 54428
rect 57039 54372 57069 54428
rect 56953 54348 57069 54372
rect 56953 54292 56983 54348
rect 57039 54292 57069 54348
rect 56953 54264 57069 54292
rect 57795 54588 57911 54616
rect 57795 54532 57825 54588
rect 57881 54532 57911 54588
rect 57795 54508 57911 54532
rect 57795 54452 57825 54508
rect 57881 54452 57911 54508
rect 57795 54428 57911 54452
rect 57795 54372 57825 54428
rect 57881 54372 57911 54428
rect 57795 54348 57911 54372
rect 57795 54292 57825 54348
rect 57881 54292 57911 54348
rect 57795 54264 57911 54292
rect 58461 54588 58525 54616
rect 58461 54532 58465 54588
rect 58521 54532 58525 54588
rect 58461 54508 58525 54532
rect 58461 54452 58465 54508
rect 58521 54452 58525 54508
rect 58461 54428 58525 54452
rect 58461 54372 58465 54428
rect 58521 54372 58525 54428
rect 58461 54348 58525 54372
rect 58461 54292 58465 54348
rect 58521 54292 58525 54348
rect 58461 54264 58525 54292
rect 59018 54588 59134 54616
rect 59018 54532 59048 54588
rect 59104 54532 59134 54588
rect 59018 54508 59134 54532
rect 59018 54452 59048 54508
rect 59104 54452 59134 54508
rect 59018 54428 59134 54452
rect 59018 54372 59048 54428
rect 59104 54372 59134 54428
rect 59018 54348 59134 54372
rect 59018 54292 59048 54348
rect 59104 54292 59134 54348
rect 59018 54264 59134 54292
rect 60296 54588 60412 54616
rect 60296 54532 60326 54588
rect 60382 54532 60412 54588
rect 60296 54508 60412 54532
rect 60296 54452 60326 54508
rect 60382 54452 60412 54508
rect 60296 54428 60412 54452
rect 60296 54372 60326 54428
rect 60382 54372 60412 54428
rect 60296 54348 60412 54372
rect 60296 54292 60326 54348
rect 60382 54292 60412 54348
rect 60296 54264 60412 54292
rect 60454 54588 60570 54616
rect 60454 54532 60484 54588
rect 60540 54532 60570 54588
rect 60454 54508 60570 54532
rect 60454 54452 60484 54508
rect 60540 54452 60570 54508
rect 60454 54428 60570 54452
rect 60454 54372 60484 54428
rect 60540 54372 60570 54428
rect 60454 54348 60570 54372
rect 60454 54292 60484 54348
rect 60540 54292 60570 54348
rect 60454 54264 60570 54292
rect 62509 54588 62683 54616
rect 62509 54532 62528 54588
rect 62584 54532 62608 54588
rect 62664 54532 62683 54588
rect 62509 54508 62683 54532
rect 62509 54452 62528 54508
rect 62584 54452 62608 54508
rect 62664 54452 62683 54508
rect 62509 54428 62683 54452
rect 62509 54372 62528 54428
rect 62584 54372 62608 54428
rect 62664 54372 62683 54428
rect 62509 54348 62683 54372
rect 62509 54292 62528 54348
rect 62584 54292 62608 54348
rect 62664 54292 62683 54348
rect 62509 54264 62683 54292
rect 2152 52236 2352 52264
rect 2152 52180 2184 52236
rect 2240 52180 2264 52236
rect 2320 52180 2352 52236
rect 2152 52156 2352 52180
rect 2152 52100 2184 52156
rect 2240 52100 2264 52156
rect 2320 52100 2352 52156
rect 2152 52076 2352 52100
rect 2152 52020 2184 52076
rect 2240 52020 2264 52076
rect 2320 52020 2352 52076
rect 2152 51996 2352 52020
rect 2152 51940 2184 51996
rect 2240 51940 2264 51996
rect 2320 51940 2352 51996
rect 2152 51912 2352 51940
rect 5374 52236 5468 52264
rect 5374 52180 5393 52236
rect 5449 52180 5468 52236
rect 5374 52156 5468 52180
rect 5374 52100 5393 52156
rect 5449 52100 5468 52156
rect 5374 52076 5468 52100
rect 5374 52020 5393 52076
rect 5449 52020 5468 52076
rect 5374 51996 5468 52020
rect 5374 51940 5393 51996
rect 5449 51940 5468 51996
rect 5374 51912 5468 51940
rect 8264 52236 8358 52264
rect 8264 52180 8283 52236
rect 8339 52180 8358 52236
rect 8264 52156 8358 52180
rect 8264 52100 8283 52156
rect 8339 52100 8358 52156
rect 8264 52076 8358 52100
rect 8264 52020 8283 52076
rect 8339 52020 8358 52076
rect 8264 51996 8358 52020
rect 8264 51940 8283 51996
rect 8339 51940 8358 51996
rect 8264 51912 8358 51940
rect 11154 52236 11248 52264
rect 11154 52180 11173 52236
rect 11229 52180 11248 52236
rect 11154 52156 11248 52180
rect 11154 52100 11173 52156
rect 11229 52100 11248 52156
rect 11154 52076 11248 52100
rect 11154 52020 11173 52076
rect 11229 52020 11248 52076
rect 11154 51996 11248 52020
rect 11154 51940 11173 51996
rect 11229 51940 11248 51996
rect 11154 51912 11248 51940
rect 14044 52236 14138 52264
rect 14044 52180 14063 52236
rect 14119 52180 14138 52236
rect 14044 52156 14138 52180
rect 14044 52100 14063 52156
rect 14119 52100 14138 52156
rect 14044 52076 14138 52100
rect 14044 52020 14063 52076
rect 14119 52020 14138 52076
rect 14044 51996 14138 52020
rect 14044 51940 14063 51996
rect 14119 51940 14138 51996
rect 14044 51912 14138 51940
rect 16934 52236 17028 52264
rect 16934 52180 16953 52236
rect 17009 52180 17028 52236
rect 16934 52156 17028 52180
rect 16934 52100 16953 52156
rect 17009 52100 17028 52156
rect 16934 52076 17028 52100
rect 16934 52020 16953 52076
rect 17009 52020 17028 52076
rect 16934 51996 17028 52020
rect 16934 51940 16953 51996
rect 17009 51940 17028 51996
rect 16934 51912 17028 51940
rect 19824 52236 19918 52264
rect 19824 52180 19843 52236
rect 19899 52180 19918 52236
rect 19824 52156 19918 52180
rect 19824 52100 19843 52156
rect 19899 52100 19918 52156
rect 19824 52076 19918 52100
rect 19824 52020 19843 52076
rect 19899 52020 19918 52076
rect 19824 51996 19918 52020
rect 19824 51940 19843 51996
rect 19899 51940 19918 51996
rect 19824 51912 19918 51940
rect 22714 52236 22808 52264
rect 22714 52180 22733 52236
rect 22789 52180 22808 52236
rect 22714 52156 22808 52180
rect 22714 52100 22733 52156
rect 22789 52100 22808 52156
rect 22714 52076 22808 52100
rect 22714 52020 22733 52076
rect 22789 52020 22808 52076
rect 22714 51996 22808 52020
rect 22714 51940 22733 51996
rect 22789 51940 22808 51996
rect 22714 51912 22808 51940
rect 25604 52236 25698 52264
rect 25604 52180 25623 52236
rect 25679 52180 25698 52236
rect 25604 52156 25698 52180
rect 25604 52100 25623 52156
rect 25679 52100 25698 52156
rect 25604 52076 25698 52100
rect 25604 52020 25623 52076
rect 25679 52020 25698 52076
rect 25604 51996 25698 52020
rect 25604 51940 25623 51996
rect 25679 51940 25698 51996
rect 25604 51912 25698 51940
rect 28494 52236 28588 52264
rect 28494 52180 28513 52236
rect 28569 52180 28588 52236
rect 28494 52156 28588 52180
rect 28494 52100 28513 52156
rect 28569 52100 28588 52156
rect 28494 52076 28588 52100
rect 28494 52020 28513 52076
rect 28569 52020 28588 52076
rect 28494 51996 28588 52020
rect 28494 51940 28513 51996
rect 28569 51940 28588 51996
rect 28494 51912 28588 51940
rect 31384 52236 31478 52264
rect 31384 52180 31403 52236
rect 31459 52180 31478 52236
rect 31384 52156 31478 52180
rect 31384 52100 31403 52156
rect 31459 52100 31478 52156
rect 31384 52076 31478 52100
rect 31384 52020 31403 52076
rect 31459 52020 31478 52076
rect 31384 51996 31478 52020
rect 31384 51940 31403 51996
rect 31459 51940 31478 51996
rect 31384 51912 31478 51940
rect 34274 52236 34368 52264
rect 34274 52180 34293 52236
rect 34349 52180 34368 52236
rect 34274 52156 34368 52180
rect 34274 52100 34293 52156
rect 34349 52100 34368 52156
rect 34274 52076 34368 52100
rect 34274 52020 34293 52076
rect 34349 52020 34368 52076
rect 34274 51996 34368 52020
rect 34274 51940 34293 51996
rect 34349 51940 34368 51996
rect 34274 51912 34368 51940
rect 37164 52236 37258 52264
rect 37164 52180 37183 52236
rect 37239 52180 37258 52236
rect 37164 52156 37258 52180
rect 37164 52100 37183 52156
rect 37239 52100 37258 52156
rect 37164 52076 37258 52100
rect 37164 52020 37183 52076
rect 37239 52020 37258 52076
rect 37164 51996 37258 52020
rect 37164 51940 37183 51996
rect 37239 51940 37258 51996
rect 37164 51912 37258 51940
rect 40054 52236 40148 52264
rect 40054 52180 40073 52236
rect 40129 52180 40148 52236
rect 40054 52156 40148 52180
rect 40054 52100 40073 52156
rect 40129 52100 40148 52156
rect 40054 52076 40148 52100
rect 40054 52020 40073 52076
rect 40129 52020 40148 52076
rect 40054 51996 40148 52020
rect 40054 51940 40073 51996
rect 40129 51940 40148 51996
rect 40054 51912 40148 51940
rect 42944 52236 43038 52264
rect 42944 52180 42963 52236
rect 43019 52180 43038 52236
rect 42944 52156 43038 52180
rect 42944 52100 42963 52156
rect 43019 52100 43038 52156
rect 42944 52076 43038 52100
rect 42944 52020 42963 52076
rect 43019 52020 43038 52076
rect 42944 51996 43038 52020
rect 42944 51940 42963 51996
rect 43019 51940 43038 51996
rect 42944 51912 43038 51940
rect 45834 52236 45928 52264
rect 45834 52180 45853 52236
rect 45909 52180 45928 52236
rect 45834 52156 45928 52180
rect 45834 52100 45853 52156
rect 45909 52100 45928 52156
rect 45834 52076 45928 52100
rect 45834 52020 45853 52076
rect 45909 52020 45928 52076
rect 45834 51996 45928 52020
rect 45834 51940 45853 51996
rect 45909 51940 45928 51996
rect 45834 51912 45928 51940
rect 48781 52236 48875 52264
rect 48781 52180 48800 52236
rect 48856 52180 48875 52236
rect 48781 52156 48875 52180
rect 48781 52100 48800 52156
rect 48856 52100 48875 52156
rect 48781 52076 48875 52100
rect 48781 52020 48800 52076
rect 48856 52020 48875 52076
rect 48781 51996 48875 52020
rect 48781 51940 48800 51996
rect 48856 51940 48875 51996
rect 48781 51912 48875 51940
rect 49630 52236 49830 52264
rect 49630 52180 49662 52236
rect 49718 52180 49742 52236
rect 49798 52180 49830 52236
rect 49630 52156 49830 52180
rect 49630 52100 49662 52156
rect 49718 52100 49742 52156
rect 49798 52100 49830 52156
rect 49630 52076 49830 52100
rect 49630 52020 49662 52076
rect 49718 52020 49742 52076
rect 49798 52020 49830 52076
rect 49630 51996 49830 52020
rect 49630 51940 49662 51996
rect 49718 51940 49742 51996
rect 49798 51940 49830 51996
rect 49630 51912 49830 51940
rect 52920 52236 53048 52264
rect 52920 52180 52956 52236
rect 53012 52180 53048 52236
rect 52920 52156 53048 52180
rect 52920 52100 52956 52156
rect 53012 52100 53048 52156
rect 52920 52076 53048 52100
rect 52920 52020 52956 52076
rect 53012 52020 53048 52076
rect 52920 51996 53048 52020
rect 52920 51940 52956 51996
rect 53012 51940 53048 51996
rect 52920 51912 53048 51940
rect 53078 52236 53206 52264
rect 53078 52180 53114 52236
rect 53170 52180 53206 52236
rect 53078 52156 53206 52180
rect 53078 52100 53114 52156
rect 53170 52100 53206 52156
rect 53078 52076 53206 52100
rect 53078 52020 53114 52076
rect 53170 52020 53206 52076
rect 53078 51996 53206 52020
rect 53078 51940 53114 51996
rect 53170 51940 53206 51996
rect 53078 51912 53206 51940
rect 53434 52236 53562 52264
rect 53434 52180 53470 52236
rect 53526 52180 53562 52236
rect 53434 52156 53562 52180
rect 53434 52100 53470 52156
rect 53526 52100 53562 52156
rect 53434 52076 53562 52100
rect 53434 52020 53470 52076
rect 53526 52020 53562 52076
rect 53434 51996 53562 52020
rect 53434 51940 53470 51996
rect 53526 51940 53562 51996
rect 53434 51912 53562 51940
rect 54752 52236 54880 52264
rect 54752 52180 54788 52236
rect 54844 52180 54880 52236
rect 54752 52156 54880 52180
rect 54752 52100 54788 52156
rect 54844 52100 54880 52156
rect 54752 52076 54880 52100
rect 54752 52020 54788 52076
rect 54844 52020 54880 52076
rect 54752 51996 54880 52020
rect 54752 51940 54788 51996
rect 54844 51940 54880 51996
rect 54752 51912 54880 51940
rect 55345 52236 55473 52264
rect 55345 52180 55381 52236
rect 55437 52180 55473 52236
rect 55345 52156 55473 52180
rect 55345 52100 55381 52156
rect 55437 52100 55473 52156
rect 55345 52076 55473 52100
rect 55345 52020 55381 52076
rect 55437 52020 55473 52076
rect 55345 51996 55473 52020
rect 55345 51940 55381 51996
rect 55437 51940 55473 51996
rect 55345 51912 55473 51940
rect 56491 52236 56619 52264
rect 56491 52180 56527 52236
rect 56583 52180 56619 52236
rect 56491 52156 56619 52180
rect 56491 52100 56527 52156
rect 56583 52100 56619 52156
rect 56491 52076 56619 52100
rect 56491 52020 56527 52076
rect 56583 52020 56619 52076
rect 56491 51996 56619 52020
rect 56491 51940 56527 51996
rect 56583 51940 56619 51996
rect 56491 51912 56619 51940
rect 57941 52236 58121 52264
rect 57941 52180 57963 52236
rect 58019 52180 58043 52236
rect 58099 52180 58121 52236
rect 57941 52156 58121 52180
rect 57941 52100 57963 52156
rect 58019 52100 58043 52156
rect 58099 52100 58121 52156
rect 57941 52076 58121 52100
rect 57941 52020 57963 52076
rect 58019 52020 58043 52076
rect 58099 52020 58121 52076
rect 57941 51996 58121 52020
rect 57941 51940 57963 51996
rect 58019 51940 58043 51996
rect 58099 51940 58121 51996
rect 57941 51912 58121 51940
rect 59164 52236 59304 52264
rect 59164 52180 59206 52236
rect 59262 52180 59304 52236
rect 59164 52156 59304 52180
rect 59164 52100 59206 52156
rect 59262 52100 59304 52156
rect 59164 52076 59304 52100
rect 59164 52020 59206 52076
rect 59262 52020 59304 52076
rect 59164 51996 59304 52020
rect 59164 51940 59206 51996
rect 59262 51940 59304 51996
rect 59164 51912 59304 51940
rect 59334 52236 59450 52264
rect 59334 52180 59364 52236
rect 59420 52180 59450 52236
rect 59334 52156 59450 52180
rect 59334 52100 59364 52156
rect 59420 52100 59450 52156
rect 59334 52076 59450 52100
rect 59334 52020 59364 52076
rect 59420 52020 59450 52076
rect 59334 51996 59450 52020
rect 59334 51940 59364 51996
rect 59420 51940 59450 51996
rect 59334 51912 59450 51940
rect 59642 52236 59758 52264
rect 59642 52180 59672 52236
rect 59728 52180 59758 52236
rect 59642 52156 59758 52180
rect 59642 52100 59672 52156
rect 59728 52100 59758 52156
rect 59642 52076 59758 52100
rect 59642 52020 59672 52076
rect 59728 52020 59758 52076
rect 59642 51996 59758 52020
rect 59642 51940 59672 51996
rect 59728 51940 59758 51996
rect 59642 51912 59758 51940
rect 59788 52236 59904 52264
rect 59788 52180 59818 52236
rect 59874 52180 59904 52236
rect 59788 52156 59904 52180
rect 59788 52100 59818 52156
rect 59874 52100 59904 52156
rect 59788 52076 59904 52100
rect 59788 52020 59818 52076
rect 59874 52020 59904 52076
rect 59788 51996 59904 52020
rect 59788 51940 59818 51996
rect 59874 51940 59904 51996
rect 59788 51912 59904 51940
rect 59934 52236 60110 52264
rect 59934 52180 59954 52236
rect 60010 52180 60034 52236
rect 60090 52180 60110 52236
rect 59934 52156 60110 52180
rect 59934 52100 59954 52156
rect 60010 52100 60034 52156
rect 60090 52100 60110 52156
rect 59934 52076 60110 52100
rect 59934 52020 59954 52076
rect 60010 52020 60034 52076
rect 60090 52020 60110 52076
rect 59934 51996 60110 52020
rect 59934 51940 59954 51996
rect 60010 51940 60034 51996
rect 60090 51940 60110 51996
rect 59934 51912 60110 51940
rect 62307 52236 62481 52264
rect 62307 52180 62326 52236
rect 62382 52180 62406 52236
rect 62462 52180 62481 52236
rect 62307 52156 62481 52180
rect 62307 52100 62326 52156
rect 62382 52100 62406 52156
rect 62462 52100 62481 52156
rect 62307 52076 62481 52100
rect 62307 52020 62326 52076
rect 62382 52020 62406 52076
rect 62462 52020 62481 52076
rect 62307 51996 62481 52020
rect 62307 51940 62326 51996
rect 62382 51940 62406 51996
rect 62462 51940 62481 51996
rect 62307 51912 62481 51940
rect 63408 49224 63460 49230
rect 63408 49166 63460 49172
rect 63420 48747 63448 49166
rect 63408 48741 63460 48747
rect 63408 48683 63460 48689
rect 63408 47325 63460 47331
rect 63408 47267 63460 47273
rect 2020 44588 2124 44616
rect 2020 44532 2044 44588
rect 2100 44532 2124 44588
rect 2020 44508 2124 44532
rect 2020 44452 2044 44508
rect 2100 44452 2124 44508
rect 2020 44428 2124 44452
rect 2020 44372 2044 44428
rect 2100 44372 2124 44428
rect 2020 44348 2124 44372
rect 2020 44292 2044 44348
rect 2100 44292 2124 44348
rect 2020 44264 2124 44292
rect 5521 44588 5615 44616
rect 5521 44532 5540 44588
rect 5596 44532 5615 44588
rect 5521 44508 5615 44532
rect 5521 44452 5540 44508
rect 5596 44452 5615 44508
rect 5521 44428 5615 44452
rect 5521 44372 5540 44428
rect 5596 44372 5615 44428
rect 5521 44348 5615 44372
rect 5521 44292 5540 44348
rect 5596 44292 5615 44348
rect 5521 44264 5615 44292
rect 8411 44588 8505 44616
rect 8411 44532 8430 44588
rect 8486 44532 8505 44588
rect 8411 44508 8505 44532
rect 8411 44452 8430 44508
rect 8486 44452 8505 44508
rect 8411 44428 8505 44452
rect 8411 44372 8430 44428
rect 8486 44372 8505 44428
rect 8411 44348 8505 44372
rect 8411 44292 8430 44348
rect 8486 44292 8505 44348
rect 8411 44264 8505 44292
rect 11301 44588 11395 44616
rect 11301 44532 11320 44588
rect 11376 44532 11395 44588
rect 11301 44508 11395 44532
rect 11301 44452 11320 44508
rect 11376 44452 11395 44508
rect 11301 44428 11395 44452
rect 11301 44372 11320 44428
rect 11376 44372 11395 44428
rect 11301 44348 11395 44372
rect 11301 44292 11320 44348
rect 11376 44292 11395 44348
rect 11301 44264 11395 44292
rect 14191 44588 14285 44616
rect 14191 44532 14210 44588
rect 14266 44532 14285 44588
rect 14191 44508 14285 44532
rect 14191 44452 14210 44508
rect 14266 44452 14285 44508
rect 14191 44428 14285 44452
rect 14191 44372 14210 44428
rect 14266 44372 14285 44428
rect 14191 44348 14285 44372
rect 14191 44292 14210 44348
rect 14266 44292 14285 44348
rect 14191 44264 14285 44292
rect 17081 44588 17175 44616
rect 17081 44532 17100 44588
rect 17156 44532 17175 44588
rect 17081 44508 17175 44532
rect 17081 44452 17100 44508
rect 17156 44452 17175 44508
rect 17081 44428 17175 44452
rect 17081 44372 17100 44428
rect 17156 44372 17175 44428
rect 17081 44348 17175 44372
rect 17081 44292 17100 44348
rect 17156 44292 17175 44348
rect 17081 44264 17175 44292
rect 19971 44588 20065 44616
rect 19971 44532 19990 44588
rect 20046 44532 20065 44588
rect 19971 44508 20065 44532
rect 19971 44452 19990 44508
rect 20046 44452 20065 44508
rect 19971 44428 20065 44452
rect 19971 44372 19990 44428
rect 20046 44372 20065 44428
rect 19971 44348 20065 44372
rect 19971 44292 19990 44348
rect 20046 44292 20065 44348
rect 19971 44264 20065 44292
rect 22861 44588 22955 44616
rect 22861 44532 22880 44588
rect 22936 44532 22955 44588
rect 22861 44508 22955 44532
rect 22861 44452 22880 44508
rect 22936 44452 22955 44508
rect 22861 44428 22955 44452
rect 22861 44372 22880 44428
rect 22936 44372 22955 44428
rect 22861 44348 22955 44372
rect 22861 44292 22880 44348
rect 22936 44292 22955 44348
rect 22861 44264 22955 44292
rect 25751 44588 25845 44616
rect 25751 44532 25770 44588
rect 25826 44532 25845 44588
rect 25751 44508 25845 44532
rect 25751 44452 25770 44508
rect 25826 44452 25845 44508
rect 25751 44428 25845 44452
rect 25751 44372 25770 44428
rect 25826 44372 25845 44428
rect 25751 44348 25845 44372
rect 25751 44292 25770 44348
rect 25826 44292 25845 44348
rect 25751 44264 25845 44292
rect 28641 44588 28735 44616
rect 28641 44532 28660 44588
rect 28716 44532 28735 44588
rect 28641 44508 28735 44532
rect 28641 44452 28660 44508
rect 28716 44452 28735 44508
rect 28641 44428 28735 44452
rect 28641 44372 28660 44428
rect 28716 44372 28735 44428
rect 28641 44348 28735 44372
rect 28641 44292 28660 44348
rect 28716 44292 28735 44348
rect 28641 44264 28735 44292
rect 31531 44588 31625 44616
rect 31531 44532 31550 44588
rect 31606 44532 31625 44588
rect 31531 44508 31625 44532
rect 31531 44452 31550 44508
rect 31606 44452 31625 44508
rect 31531 44428 31625 44452
rect 31531 44372 31550 44428
rect 31606 44372 31625 44428
rect 31531 44348 31625 44372
rect 31531 44292 31550 44348
rect 31606 44292 31625 44348
rect 31531 44264 31625 44292
rect 34421 44588 34515 44616
rect 34421 44532 34440 44588
rect 34496 44532 34515 44588
rect 34421 44508 34515 44532
rect 34421 44452 34440 44508
rect 34496 44452 34515 44508
rect 34421 44428 34515 44452
rect 34421 44372 34440 44428
rect 34496 44372 34515 44428
rect 34421 44348 34515 44372
rect 34421 44292 34440 44348
rect 34496 44292 34515 44348
rect 34421 44264 34515 44292
rect 37311 44588 37405 44616
rect 37311 44532 37330 44588
rect 37386 44532 37405 44588
rect 37311 44508 37405 44532
rect 37311 44452 37330 44508
rect 37386 44452 37405 44508
rect 37311 44428 37405 44452
rect 37311 44372 37330 44428
rect 37386 44372 37405 44428
rect 37311 44348 37405 44372
rect 37311 44292 37330 44348
rect 37386 44292 37405 44348
rect 37311 44264 37405 44292
rect 40201 44588 40295 44616
rect 40201 44532 40220 44588
rect 40276 44532 40295 44588
rect 40201 44508 40295 44532
rect 40201 44452 40220 44508
rect 40276 44452 40295 44508
rect 40201 44428 40295 44452
rect 40201 44372 40220 44428
rect 40276 44372 40295 44428
rect 40201 44348 40295 44372
rect 40201 44292 40220 44348
rect 40276 44292 40295 44348
rect 40201 44264 40295 44292
rect 43091 44588 43185 44616
rect 43091 44532 43110 44588
rect 43166 44532 43185 44588
rect 43091 44508 43185 44532
rect 43091 44452 43110 44508
rect 43166 44452 43185 44508
rect 43091 44428 43185 44452
rect 43091 44372 43110 44428
rect 43166 44372 43185 44428
rect 43091 44348 43185 44372
rect 43091 44292 43110 44348
rect 43166 44292 43185 44348
rect 43091 44264 43185 44292
rect 45981 44588 46075 44616
rect 45981 44532 46000 44588
rect 46056 44532 46075 44588
rect 45981 44508 46075 44532
rect 45981 44452 46000 44508
rect 46056 44452 46075 44508
rect 45981 44428 46075 44452
rect 45981 44372 46000 44428
rect 46056 44372 46075 44428
rect 45981 44348 46075 44372
rect 45981 44292 46000 44348
rect 46056 44292 46075 44348
rect 45981 44264 46075 44292
rect 52210 44588 52320 44616
rect 52210 44532 52237 44588
rect 52293 44532 52320 44588
rect 52210 44508 52320 44532
rect 52210 44452 52237 44508
rect 52293 44452 52320 44508
rect 52210 44428 52320 44452
rect 52210 44372 52237 44428
rect 52293 44372 52320 44428
rect 52210 44348 52320 44372
rect 52210 44292 52237 44348
rect 52293 44292 52320 44348
rect 52210 44264 52320 44292
rect 53602 44588 53730 44616
rect 53602 44532 53638 44588
rect 53694 44532 53730 44588
rect 53602 44508 53730 44532
rect 53602 44452 53638 44508
rect 53694 44452 53730 44508
rect 53602 44428 53730 44452
rect 53602 44372 53638 44428
rect 53694 44372 53730 44428
rect 53602 44348 53730 44372
rect 53602 44292 53638 44348
rect 53694 44292 53730 44348
rect 53602 44264 53730 44292
rect 54514 44588 54642 44616
rect 54514 44532 54550 44588
rect 54606 44532 54642 44588
rect 54514 44508 54642 44532
rect 54514 44452 54550 44508
rect 54606 44452 54642 44508
rect 54514 44428 54642 44452
rect 54514 44372 54550 44428
rect 54606 44372 54642 44428
rect 54514 44348 54642 44372
rect 54514 44292 54550 44348
rect 54606 44292 54642 44348
rect 54514 44264 54642 44292
rect 54910 44588 55026 44616
rect 54910 44532 54940 44588
rect 54996 44532 55026 44588
rect 54910 44508 55026 44532
rect 54910 44452 54940 44508
rect 54996 44452 55026 44508
rect 54910 44428 55026 44452
rect 54910 44372 54940 44428
rect 54996 44372 55026 44428
rect 54910 44348 55026 44372
rect 54910 44292 54940 44348
rect 54996 44292 55026 44348
rect 54910 44264 55026 44292
rect 55620 44588 55748 44616
rect 55620 44532 55656 44588
rect 55712 44532 55748 44588
rect 55620 44508 55748 44532
rect 55620 44452 55656 44508
rect 55712 44452 55748 44508
rect 55620 44428 55748 44452
rect 55620 44372 55656 44428
rect 55712 44372 55748 44428
rect 55620 44348 55748 44372
rect 55620 44292 55656 44348
rect 55712 44292 55748 44348
rect 55620 44264 55748 44292
rect 56198 44588 56326 44616
rect 56198 44532 56234 44588
rect 56290 44532 56326 44588
rect 56198 44508 56326 44532
rect 56198 44452 56234 44508
rect 56290 44452 56326 44508
rect 56198 44428 56326 44452
rect 56198 44372 56234 44428
rect 56290 44372 56326 44428
rect 56198 44348 56326 44372
rect 56198 44292 56234 44348
rect 56290 44292 56326 44348
rect 56198 44264 56326 44292
rect 56649 44588 56765 44616
rect 56649 44532 56679 44588
rect 56735 44532 56765 44588
rect 56649 44508 56765 44532
rect 56649 44452 56679 44508
rect 56735 44452 56765 44508
rect 56649 44428 56765 44452
rect 56649 44372 56679 44428
rect 56735 44372 56765 44428
rect 56649 44348 56765 44372
rect 56649 44292 56679 44348
rect 56735 44292 56765 44348
rect 56649 44264 56765 44292
rect 56953 44588 57069 44616
rect 56953 44532 56983 44588
rect 57039 44532 57069 44588
rect 56953 44508 57069 44532
rect 56953 44452 56983 44508
rect 57039 44452 57069 44508
rect 56953 44428 57069 44452
rect 56953 44372 56983 44428
rect 57039 44372 57069 44428
rect 56953 44348 57069 44372
rect 56953 44292 56983 44348
rect 57039 44292 57069 44348
rect 56953 44264 57069 44292
rect 57795 44588 57911 44616
rect 57795 44532 57825 44588
rect 57881 44532 57911 44588
rect 57795 44508 57911 44532
rect 57795 44452 57825 44508
rect 57881 44452 57911 44508
rect 57795 44428 57911 44452
rect 57795 44372 57825 44428
rect 57881 44372 57911 44428
rect 57795 44348 57911 44372
rect 57795 44292 57825 44348
rect 57881 44292 57911 44348
rect 57795 44264 57911 44292
rect 58345 44588 58409 44616
rect 58345 44532 58349 44588
rect 58405 44532 58409 44588
rect 58345 44508 58409 44532
rect 58345 44452 58349 44508
rect 58405 44452 58409 44508
rect 58345 44428 58409 44452
rect 58345 44372 58349 44428
rect 58405 44372 58409 44428
rect 58345 44348 58409 44372
rect 58345 44292 58349 44348
rect 58405 44292 58409 44348
rect 58345 44264 58409 44292
rect 59018 44588 59134 44616
rect 59018 44532 59048 44588
rect 59104 44532 59134 44588
rect 59018 44508 59134 44532
rect 59018 44452 59048 44508
rect 59104 44452 59134 44508
rect 59018 44428 59134 44452
rect 59018 44372 59048 44428
rect 59104 44372 59134 44428
rect 59018 44348 59134 44372
rect 59018 44292 59048 44348
rect 59104 44292 59134 44348
rect 59018 44264 59134 44292
rect 60296 44588 60412 44616
rect 60296 44532 60326 44588
rect 60382 44532 60412 44588
rect 60296 44508 60412 44532
rect 60296 44452 60326 44508
rect 60382 44452 60412 44508
rect 60296 44428 60412 44452
rect 60296 44372 60326 44428
rect 60382 44372 60412 44428
rect 60296 44348 60412 44372
rect 60296 44292 60326 44348
rect 60382 44292 60412 44348
rect 60296 44264 60412 44292
rect 60454 44588 60570 44616
rect 60454 44532 60484 44588
rect 60540 44532 60570 44588
rect 60454 44508 60570 44532
rect 60454 44452 60484 44508
rect 60540 44452 60570 44508
rect 60454 44428 60570 44452
rect 60454 44372 60484 44428
rect 60540 44372 60570 44428
rect 60454 44348 60570 44372
rect 60454 44292 60484 44348
rect 60540 44292 60570 44348
rect 60454 44264 60570 44292
rect 62509 44588 62683 44616
rect 62509 44532 62528 44588
rect 62584 44532 62608 44588
rect 62664 44532 62683 44588
rect 62509 44508 62683 44532
rect 62509 44452 62528 44508
rect 62584 44452 62608 44508
rect 62664 44452 62683 44508
rect 62509 44428 62683 44452
rect 62509 44372 62528 44428
rect 62584 44372 62608 44428
rect 62664 44372 62683 44428
rect 62509 44348 62683 44372
rect 62509 44292 62528 44348
rect 62584 44292 62608 44348
rect 62664 44292 62683 44348
rect 62509 44264 62683 44292
rect 2152 42236 2352 42264
rect 2152 42180 2184 42236
rect 2240 42180 2264 42236
rect 2320 42180 2352 42236
rect 2152 42156 2352 42180
rect 2152 42100 2184 42156
rect 2240 42100 2264 42156
rect 2320 42100 2352 42156
rect 2152 42076 2352 42100
rect 2152 42020 2184 42076
rect 2240 42020 2264 42076
rect 2320 42020 2352 42076
rect 2152 41996 2352 42020
rect 2152 41940 2184 41996
rect 2240 41940 2264 41996
rect 2320 41940 2352 41996
rect 2152 41912 2352 41940
rect 5374 42236 5468 42264
rect 5374 42180 5393 42236
rect 5449 42180 5468 42236
rect 5374 42156 5468 42180
rect 5374 42100 5393 42156
rect 5449 42100 5468 42156
rect 5374 42076 5468 42100
rect 5374 42020 5393 42076
rect 5449 42020 5468 42076
rect 5374 41996 5468 42020
rect 5374 41940 5393 41996
rect 5449 41940 5468 41996
rect 5374 41912 5468 41940
rect 8264 42236 8358 42264
rect 8264 42180 8283 42236
rect 8339 42180 8358 42236
rect 8264 42156 8358 42180
rect 8264 42100 8283 42156
rect 8339 42100 8358 42156
rect 8264 42076 8358 42100
rect 8264 42020 8283 42076
rect 8339 42020 8358 42076
rect 8264 41996 8358 42020
rect 8264 41940 8283 41996
rect 8339 41940 8358 41996
rect 8264 41912 8358 41940
rect 11154 42236 11248 42264
rect 11154 42180 11173 42236
rect 11229 42180 11248 42236
rect 11154 42156 11248 42180
rect 11154 42100 11173 42156
rect 11229 42100 11248 42156
rect 11154 42076 11248 42100
rect 11154 42020 11173 42076
rect 11229 42020 11248 42076
rect 11154 41996 11248 42020
rect 11154 41940 11173 41996
rect 11229 41940 11248 41996
rect 11154 41912 11248 41940
rect 14044 42236 14138 42264
rect 14044 42180 14063 42236
rect 14119 42180 14138 42236
rect 14044 42156 14138 42180
rect 14044 42100 14063 42156
rect 14119 42100 14138 42156
rect 14044 42076 14138 42100
rect 14044 42020 14063 42076
rect 14119 42020 14138 42076
rect 14044 41996 14138 42020
rect 14044 41940 14063 41996
rect 14119 41940 14138 41996
rect 14044 41912 14138 41940
rect 16934 42236 17028 42264
rect 16934 42180 16953 42236
rect 17009 42180 17028 42236
rect 16934 42156 17028 42180
rect 16934 42100 16953 42156
rect 17009 42100 17028 42156
rect 16934 42076 17028 42100
rect 16934 42020 16953 42076
rect 17009 42020 17028 42076
rect 16934 41996 17028 42020
rect 16934 41940 16953 41996
rect 17009 41940 17028 41996
rect 16934 41912 17028 41940
rect 19824 42236 19918 42264
rect 19824 42180 19843 42236
rect 19899 42180 19918 42236
rect 19824 42156 19918 42180
rect 19824 42100 19843 42156
rect 19899 42100 19918 42156
rect 19824 42076 19918 42100
rect 19824 42020 19843 42076
rect 19899 42020 19918 42076
rect 19824 41996 19918 42020
rect 19824 41940 19843 41996
rect 19899 41940 19918 41996
rect 19824 41912 19918 41940
rect 22714 42236 22808 42264
rect 22714 42180 22733 42236
rect 22789 42180 22808 42236
rect 22714 42156 22808 42180
rect 22714 42100 22733 42156
rect 22789 42100 22808 42156
rect 22714 42076 22808 42100
rect 22714 42020 22733 42076
rect 22789 42020 22808 42076
rect 22714 41996 22808 42020
rect 22714 41940 22733 41996
rect 22789 41940 22808 41996
rect 22714 41912 22808 41940
rect 25604 42236 25698 42264
rect 25604 42180 25623 42236
rect 25679 42180 25698 42236
rect 25604 42156 25698 42180
rect 25604 42100 25623 42156
rect 25679 42100 25698 42156
rect 25604 42076 25698 42100
rect 25604 42020 25623 42076
rect 25679 42020 25698 42076
rect 25604 41996 25698 42020
rect 25604 41940 25623 41996
rect 25679 41940 25698 41996
rect 25604 41912 25698 41940
rect 28494 42236 28588 42264
rect 28494 42180 28513 42236
rect 28569 42180 28588 42236
rect 28494 42156 28588 42180
rect 28494 42100 28513 42156
rect 28569 42100 28588 42156
rect 28494 42076 28588 42100
rect 28494 42020 28513 42076
rect 28569 42020 28588 42076
rect 28494 41996 28588 42020
rect 28494 41940 28513 41996
rect 28569 41940 28588 41996
rect 28494 41912 28588 41940
rect 31384 42236 31478 42264
rect 31384 42180 31403 42236
rect 31459 42180 31478 42236
rect 31384 42156 31478 42180
rect 31384 42100 31403 42156
rect 31459 42100 31478 42156
rect 31384 42076 31478 42100
rect 31384 42020 31403 42076
rect 31459 42020 31478 42076
rect 31384 41996 31478 42020
rect 31384 41940 31403 41996
rect 31459 41940 31478 41996
rect 31384 41912 31478 41940
rect 34274 42236 34368 42264
rect 34274 42180 34293 42236
rect 34349 42180 34368 42236
rect 34274 42156 34368 42180
rect 34274 42100 34293 42156
rect 34349 42100 34368 42156
rect 34274 42076 34368 42100
rect 34274 42020 34293 42076
rect 34349 42020 34368 42076
rect 34274 41996 34368 42020
rect 34274 41940 34293 41996
rect 34349 41940 34368 41996
rect 34274 41912 34368 41940
rect 37164 42236 37258 42264
rect 37164 42180 37183 42236
rect 37239 42180 37258 42236
rect 37164 42156 37258 42180
rect 37164 42100 37183 42156
rect 37239 42100 37258 42156
rect 37164 42076 37258 42100
rect 37164 42020 37183 42076
rect 37239 42020 37258 42076
rect 37164 41996 37258 42020
rect 37164 41940 37183 41996
rect 37239 41940 37258 41996
rect 37164 41912 37258 41940
rect 40054 42236 40148 42264
rect 40054 42180 40073 42236
rect 40129 42180 40148 42236
rect 40054 42156 40148 42180
rect 40054 42100 40073 42156
rect 40129 42100 40148 42156
rect 40054 42076 40148 42100
rect 40054 42020 40073 42076
rect 40129 42020 40148 42076
rect 40054 41996 40148 42020
rect 40054 41940 40073 41996
rect 40129 41940 40148 41996
rect 40054 41912 40148 41940
rect 42944 42236 43038 42264
rect 42944 42180 42963 42236
rect 43019 42180 43038 42236
rect 42944 42156 43038 42180
rect 42944 42100 42963 42156
rect 43019 42100 43038 42156
rect 42944 42076 43038 42100
rect 42944 42020 42963 42076
rect 43019 42020 43038 42076
rect 42944 41996 43038 42020
rect 42944 41940 42963 41996
rect 43019 41940 43038 41996
rect 42944 41912 43038 41940
rect 45834 42236 45928 42264
rect 45834 42180 45853 42236
rect 45909 42180 45928 42236
rect 45834 42156 45928 42180
rect 45834 42100 45853 42156
rect 45909 42100 45928 42156
rect 45834 42076 45928 42100
rect 45834 42020 45853 42076
rect 45909 42020 45928 42076
rect 45834 41996 45928 42020
rect 45834 41940 45853 41996
rect 45909 41940 45928 41996
rect 45834 41912 45928 41940
rect 48781 42236 48875 42264
rect 48781 42180 48800 42236
rect 48856 42180 48875 42236
rect 48781 42156 48875 42180
rect 48781 42100 48800 42156
rect 48856 42100 48875 42156
rect 48781 42076 48875 42100
rect 48781 42020 48800 42076
rect 48856 42020 48875 42076
rect 48781 41996 48875 42020
rect 48781 41940 48800 41996
rect 48856 41940 48875 41996
rect 48781 41912 48875 41940
rect 49630 42236 49830 42264
rect 49630 42180 49662 42236
rect 49718 42180 49742 42236
rect 49798 42180 49830 42236
rect 49630 42156 49830 42180
rect 49630 42100 49662 42156
rect 49718 42100 49742 42156
rect 49798 42100 49830 42156
rect 49630 42076 49830 42100
rect 49630 42020 49662 42076
rect 49718 42020 49742 42076
rect 49798 42020 49830 42076
rect 49630 41996 49830 42020
rect 49630 41940 49662 41996
rect 49718 41940 49742 41996
rect 49798 41940 49830 41996
rect 49630 41912 49830 41940
rect 52920 42236 53048 42264
rect 52920 42180 52956 42236
rect 53012 42180 53048 42236
rect 52920 42156 53048 42180
rect 52920 42100 52956 42156
rect 53012 42100 53048 42156
rect 52920 42076 53048 42100
rect 52920 42020 52956 42076
rect 53012 42020 53048 42076
rect 52920 41996 53048 42020
rect 52920 41940 52956 41996
rect 53012 41940 53048 41996
rect 52920 41912 53048 41940
rect 53078 42236 53206 42264
rect 53078 42180 53114 42236
rect 53170 42180 53206 42236
rect 53078 42156 53206 42180
rect 53078 42100 53114 42156
rect 53170 42100 53206 42156
rect 53078 42076 53206 42100
rect 53078 42020 53114 42076
rect 53170 42020 53206 42076
rect 53078 41996 53206 42020
rect 53078 41940 53114 41996
rect 53170 41940 53206 41996
rect 53078 41912 53206 41940
rect 53434 42236 53562 42264
rect 53434 42180 53470 42236
rect 53526 42180 53562 42236
rect 53434 42156 53562 42180
rect 53434 42100 53470 42156
rect 53526 42100 53562 42156
rect 53434 42076 53562 42100
rect 53434 42020 53470 42076
rect 53526 42020 53562 42076
rect 53434 41996 53562 42020
rect 53434 41940 53470 41996
rect 53526 41940 53562 41996
rect 53434 41912 53562 41940
rect 54752 42236 54880 42264
rect 54752 42180 54788 42236
rect 54844 42180 54880 42236
rect 54752 42156 54880 42180
rect 54752 42100 54788 42156
rect 54844 42100 54880 42156
rect 54752 42076 54880 42100
rect 54752 42020 54788 42076
rect 54844 42020 54880 42076
rect 54752 41996 54880 42020
rect 54752 41940 54788 41996
rect 54844 41940 54880 41996
rect 54752 41912 54880 41940
rect 55345 42236 55473 42264
rect 55345 42180 55381 42236
rect 55437 42180 55473 42236
rect 55345 42156 55473 42180
rect 55345 42100 55381 42156
rect 55437 42100 55473 42156
rect 55345 42076 55473 42100
rect 55345 42020 55381 42076
rect 55437 42020 55473 42076
rect 55345 41996 55473 42020
rect 55345 41940 55381 41996
rect 55437 41940 55473 41996
rect 55345 41912 55473 41940
rect 56491 42236 56619 42264
rect 56491 42180 56527 42236
rect 56583 42180 56619 42236
rect 56491 42156 56619 42180
rect 56491 42100 56527 42156
rect 56583 42100 56619 42156
rect 56491 42076 56619 42100
rect 56491 42020 56527 42076
rect 56583 42020 56619 42076
rect 56491 41996 56619 42020
rect 56491 41940 56527 41996
rect 56583 41940 56619 41996
rect 56491 41912 56619 41940
rect 57941 42236 58121 42264
rect 57941 42180 57963 42236
rect 58019 42180 58043 42236
rect 58099 42180 58121 42236
rect 57941 42156 58121 42180
rect 57941 42100 57963 42156
rect 58019 42100 58043 42156
rect 58099 42100 58121 42156
rect 57941 42076 58121 42100
rect 57941 42020 57963 42076
rect 58019 42020 58043 42076
rect 58099 42020 58121 42076
rect 57941 41996 58121 42020
rect 57941 41940 57963 41996
rect 58019 41940 58043 41996
rect 58099 41940 58121 41996
rect 57941 41912 58121 41940
rect 59164 42236 59304 42264
rect 59164 42180 59206 42236
rect 59262 42180 59304 42236
rect 59164 42156 59304 42180
rect 59164 42100 59206 42156
rect 59262 42100 59304 42156
rect 59164 42076 59304 42100
rect 59164 42020 59206 42076
rect 59262 42020 59304 42076
rect 59164 41996 59304 42020
rect 59164 41940 59206 41996
rect 59262 41940 59304 41996
rect 59164 41912 59304 41940
rect 59334 42236 59450 42264
rect 59334 42180 59364 42236
rect 59420 42180 59450 42236
rect 59334 42156 59450 42180
rect 59334 42100 59364 42156
rect 59420 42100 59450 42156
rect 59334 42076 59450 42100
rect 59334 42020 59364 42076
rect 59420 42020 59450 42076
rect 59334 41996 59450 42020
rect 59334 41940 59364 41996
rect 59420 41940 59450 41996
rect 59334 41912 59450 41940
rect 59642 42236 59758 42264
rect 59642 42180 59672 42236
rect 59728 42180 59758 42236
rect 59642 42156 59758 42180
rect 59642 42100 59672 42156
rect 59728 42100 59758 42156
rect 59642 42076 59758 42100
rect 59642 42020 59672 42076
rect 59728 42020 59758 42076
rect 59642 41996 59758 42020
rect 59642 41940 59672 41996
rect 59728 41940 59758 41996
rect 59642 41912 59758 41940
rect 59788 42236 59904 42264
rect 59788 42180 59818 42236
rect 59874 42180 59904 42236
rect 59788 42156 59904 42180
rect 59788 42100 59818 42156
rect 59874 42100 59904 42156
rect 59788 42076 59904 42100
rect 59788 42020 59818 42076
rect 59874 42020 59904 42076
rect 59788 41996 59904 42020
rect 59788 41940 59818 41996
rect 59874 41940 59904 41996
rect 59788 41912 59904 41940
rect 59934 42236 60110 42264
rect 59934 42180 59954 42236
rect 60010 42180 60034 42236
rect 60090 42180 60110 42236
rect 59934 42156 60110 42180
rect 59934 42100 59954 42156
rect 60010 42100 60034 42156
rect 60090 42100 60110 42156
rect 59934 42076 60110 42100
rect 59934 42020 59954 42076
rect 60010 42020 60034 42076
rect 60090 42020 60110 42076
rect 59934 41996 60110 42020
rect 59934 41940 59954 41996
rect 60010 41940 60034 41996
rect 60090 41940 60110 41996
rect 59934 41912 60110 41940
rect 62307 42236 62481 42264
rect 62307 42180 62326 42236
rect 62382 42180 62406 42236
rect 62462 42180 62481 42236
rect 62307 42156 62481 42180
rect 62307 42100 62326 42156
rect 62382 42100 62406 42156
rect 62462 42100 62481 42156
rect 62307 42076 62481 42100
rect 62307 42020 62326 42076
rect 62382 42020 62406 42076
rect 62462 42020 62481 42076
rect 62307 41996 62481 42020
rect 62307 41940 62326 41996
rect 62382 41940 62406 41996
rect 62462 41940 62481 41996
rect 62307 41912 62481 41940
rect 63420 39642 63448 47267
rect 63408 39636 63460 39642
rect 63408 39578 63460 39584
rect 63408 38936 63460 38942
rect 63408 38878 63460 38884
rect 2020 34588 2124 34616
rect 2020 34532 2044 34588
rect 2100 34532 2124 34588
rect 2020 34508 2124 34532
rect 2020 34452 2044 34508
rect 2100 34452 2124 34508
rect 2020 34428 2124 34452
rect 2020 34372 2044 34428
rect 2100 34372 2124 34428
rect 2020 34348 2124 34372
rect 2020 34292 2044 34348
rect 2100 34292 2124 34348
rect 2020 34264 2124 34292
rect 5521 34588 5615 34616
rect 5521 34532 5540 34588
rect 5596 34532 5615 34588
rect 5521 34508 5615 34532
rect 5521 34452 5540 34508
rect 5596 34452 5615 34508
rect 5521 34428 5615 34452
rect 5521 34372 5540 34428
rect 5596 34372 5615 34428
rect 5521 34348 5615 34372
rect 5521 34292 5540 34348
rect 5596 34292 5615 34348
rect 5521 34264 5615 34292
rect 8411 34588 8505 34616
rect 8411 34532 8430 34588
rect 8486 34532 8505 34588
rect 8411 34508 8505 34532
rect 8411 34452 8430 34508
rect 8486 34452 8505 34508
rect 8411 34428 8505 34452
rect 8411 34372 8430 34428
rect 8486 34372 8505 34428
rect 8411 34348 8505 34372
rect 8411 34292 8430 34348
rect 8486 34292 8505 34348
rect 8411 34264 8505 34292
rect 11301 34588 11395 34616
rect 11301 34532 11320 34588
rect 11376 34532 11395 34588
rect 11301 34508 11395 34532
rect 11301 34452 11320 34508
rect 11376 34452 11395 34508
rect 11301 34428 11395 34452
rect 11301 34372 11320 34428
rect 11376 34372 11395 34428
rect 11301 34348 11395 34372
rect 11301 34292 11320 34348
rect 11376 34292 11395 34348
rect 11301 34264 11395 34292
rect 14191 34588 14285 34616
rect 14191 34532 14210 34588
rect 14266 34532 14285 34588
rect 14191 34508 14285 34532
rect 14191 34452 14210 34508
rect 14266 34452 14285 34508
rect 14191 34428 14285 34452
rect 14191 34372 14210 34428
rect 14266 34372 14285 34428
rect 14191 34348 14285 34372
rect 14191 34292 14210 34348
rect 14266 34292 14285 34348
rect 14191 34264 14285 34292
rect 17081 34588 17175 34616
rect 17081 34532 17100 34588
rect 17156 34532 17175 34588
rect 17081 34508 17175 34532
rect 17081 34452 17100 34508
rect 17156 34452 17175 34508
rect 17081 34428 17175 34452
rect 17081 34372 17100 34428
rect 17156 34372 17175 34428
rect 17081 34348 17175 34372
rect 17081 34292 17100 34348
rect 17156 34292 17175 34348
rect 17081 34264 17175 34292
rect 19971 34588 20065 34616
rect 19971 34532 19990 34588
rect 20046 34532 20065 34588
rect 19971 34508 20065 34532
rect 19971 34452 19990 34508
rect 20046 34452 20065 34508
rect 19971 34428 20065 34452
rect 19971 34372 19990 34428
rect 20046 34372 20065 34428
rect 19971 34348 20065 34372
rect 19971 34292 19990 34348
rect 20046 34292 20065 34348
rect 19971 34264 20065 34292
rect 22861 34588 22955 34616
rect 22861 34532 22880 34588
rect 22936 34532 22955 34588
rect 22861 34508 22955 34532
rect 22861 34452 22880 34508
rect 22936 34452 22955 34508
rect 22861 34428 22955 34452
rect 22861 34372 22880 34428
rect 22936 34372 22955 34428
rect 22861 34348 22955 34372
rect 22861 34292 22880 34348
rect 22936 34292 22955 34348
rect 22861 34264 22955 34292
rect 25751 34588 25845 34616
rect 25751 34532 25770 34588
rect 25826 34532 25845 34588
rect 25751 34508 25845 34532
rect 25751 34452 25770 34508
rect 25826 34452 25845 34508
rect 25751 34428 25845 34452
rect 25751 34372 25770 34428
rect 25826 34372 25845 34428
rect 25751 34348 25845 34372
rect 25751 34292 25770 34348
rect 25826 34292 25845 34348
rect 25751 34264 25845 34292
rect 28641 34588 28735 34616
rect 28641 34532 28660 34588
rect 28716 34532 28735 34588
rect 28641 34508 28735 34532
rect 28641 34452 28660 34508
rect 28716 34452 28735 34508
rect 28641 34428 28735 34452
rect 28641 34372 28660 34428
rect 28716 34372 28735 34428
rect 28641 34348 28735 34372
rect 28641 34292 28660 34348
rect 28716 34292 28735 34348
rect 28641 34264 28735 34292
rect 31531 34588 31625 34616
rect 31531 34532 31550 34588
rect 31606 34532 31625 34588
rect 31531 34508 31625 34532
rect 31531 34452 31550 34508
rect 31606 34452 31625 34508
rect 31531 34428 31625 34452
rect 31531 34372 31550 34428
rect 31606 34372 31625 34428
rect 31531 34348 31625 34372
rect 31531 34292 31550 34348
rect 31606 34292 31625 34348
rect 31531 34264 31625 34292
rect 34421 34588 34515 34616
rect 34421 34532 34440 34588
rect 34496 34532 34515 34588
rect 34421 34508 34515 34532
rect 34421 34452 34440 34508
rect 34496 34452 34515 34508
rect 34421 34428 34515 34452
rect 34421 34372 34440 34428
rect 34496 34372 34515 34428
rect 34421 34348 34515 34372
rect 34421 34292 34440 34348
rect 34496 34292 34515 34348
rect 34421 34264 34515 34292
rect 37311 34588 37405 34616
rect 37311 34532 37330 34588
rect 37386 34532 37405 34588
rect 37311 34508 37405 34532
rect 37311 34452 37330 34508
rect 37386 34452 37405 34508
rect 37311 34428 37405 34452
rect 37311 34372 37330 34428
rect 37386 34372 37405 34428
rect 37311 34348 37405 34372
rect 37311 34292 37330 34348
rect 37386 34292 37405 34348
rect 37311 34264 37405 34292
rect 40201 34588 40295 34616
rect 40201 34532 40220 34588
rect 40276 34532 40295 34588
rect 40201 34508 40295 34532
rect 40201 34452 40220 34508
rect 40276 34452 40295 34508
rect 40201 34428 40295 34452
rect 40201 34372 40220 34428
rect 40276 34372 40295 34428
rect 40201 34348 40295 34372
rect 40201 34292 40220 34348
rect 40276 34292 40295 34348
rect 40201 34264 40295 34292
rect 43091 34588 43185 34616
rect 43091 34532 43110 34588
rect 43166 34532 43185 34588
rect 43091 34508 43185 34532
rect 43091 34452 43110 34508
rect 43166 34452 43185 34508
rect 43091 34428 43185 34452
rect 43091 34372 43110 34428
rect 43166 34372 43185 34428
rect 43091 34348 43185 34372
rect 43091 34292 43110 34348
rect 43166 34292 43185 34348
rect 43091 34264 43185 34292
rect 45981 34588 46075 34616
rect 45981 34532 46000 34588
rect 46056 34532 46075 34588
rect 45981 34508 46075 34532
rect 45981 34452 46000 34508
rect 46056 34452 46075 34508
rect 45981 34428 46075 34452
rect 45981 34372 46000 34428
rect 46056 34372 46075 34428
rect 45981 34348 46075 34372
rect 45981 34292 46000 34348
rect 46056 34292 46075 34348
rect 45981 34264 46075 34292
rect 48989 34588 49083 34616
rect 48989 34532 49008 34588
rect 49064 34532 49083 34588
rect 48989 34508 49083 34532
rect 48989 34452 49008 34508
rect 49064 34452 49083 34508
rect 48989 34428 49083 34452
rect 48989 34372 49008 34428
rect 49064 34372 49083 34428
rect 48989 34348 49083 34372
rect 48989 34292 49008 34348
rect 49064 34292 49083 34348
rect 48989 34264 49083 34292
rect 52210 34588 52320 34616
rect 52210 34532 52237 34588
rect 52293 34532 52320 34588
rect 52210 34508 52320 34532
rect 52210 34452 52237 34508
rect 52293 34452 52320 34508
rect 52210 34428 52320 34452
rect 52210 34372 52237 34428
rect 52293 34372 52320 34428
rect 52210 34348 52320 34372
rect 52210 34292 52237 34348
rect 52293 34292 52320 34348
rect 52210 34264 52320 34292
rect 53602 34588 53730 34616
rect 53602 34532 53638 34588
rect 53694 34532 53730 34588
rect 53602 34508 53730 34532
rect 53602 34452 53638 34508
rect 53694 34452 53730 34508
rect 53602 34428 53730 34452
rect 53602 34372 53638 34428
rect 53694 34372 53730 34428
rect 53602 34348 53730 34372
rect 53602 34292 53638 34348
rect 53694 34292 53730 34348
rect 53602 34264 53730 34292
rect 53770 34588 53898 34616
rect 53770 34532 53806 34588
rect 53862 34532 53898 34588
rect 53770 34508 53898 34532
rect 53770 34452 53806 34508
rect 53862 34452 53898 34508
rect 53770 34428 53898 34452
rect 53770 34372 53806 34428
rect 53862 34372 53898 34428
rect 53770 34348 53898 34372
rect 53770 34292 53806 34348
rect 53862 34292 53898 34348
rect 53770 34264 53898 34292
rect 54514 34588 54642 34616
rect 54514 34532 54550 34588
rect 54606 34532 54642 34588
rect 54514 34508 54642 34532
rect 54514 34452 54550 34508
rect 54606 34452 54642 34508
rect 54514 34428 54642 34452
rect 54514 34372 54550 34428
rect 54606 34372 54642 34428
rect 54514 34348 54642 34372
rect 54514 34292 54550 34348
rect 54606 34292 54642 34348
rect 54514 34264 54642 34292
rect 54910 34588 55026 34616
rect 54910 34532 54940 34588
rect 54996 34532 55026 34588
rect 54910 34508 55026 34532
rect 54910 34452 54940 34508
rect 54996 34452 55026 34508
rect 54910 34428 55026 34452
rect 54910 34372 54940 34428
rect 54996 34372 55026 34428
rect 54910 34348 55026 34372
rect 54910 34292 54940 34348
rect 54996 34292 55026 34348
rect 54910 34264 55026 34292
rect 55620 34588 55748 34616
rect 55620 34532 55656 34588
rect 55712 34532 55748 34588
rect 55620 34508 55748 34532
rect 55620 34452 55656 34508
rect 55712 34452 55748 34508
rect 55620 34428 55748 34452
rect 55620 34372 55656 34428
rect 55712 34372 55748 34428
rect 55620 34348 55748 34372
rect 55620 34292 55656 34348
rect 55712 34292 55748 34348
rect 55620 34264 55748 34292
rect 56198 34588 56326 34616
rect 56198 34532 56234 34588
rect 56290 34532 56326 34588
rect 56198 34508 56326 34532
rect 56198 34452 56234 34508
rect 56290 34452 56326 34508
rect 56198 34428 56326 34452
rect 56198 34372 56234 34428
rect 56290 34372 56326 34428
rect 56198 34348 56326 34372
rect 56198 34292 56234 34348
rect 56290 34292 56326 34348
rect 56198 34264 56326 34292
rect 56649 34588 56765 34616
rect 56649 34532 56679 34588
rect 56735 34532 56765 34588
rect 56649 34508 56765 34532
rect 56649 34452 56679 34508
rect 56735 34452 56765 34508
rect 56649 34428 56765 34452
rect 56649 34372 56679 34428
rect 56735 34372 56765 34428
rect 56649 34348 56765 34372
rect 56649 34292 56679 34348
rect 56735 34292 56765 34348
rect 56649 34264 56765 34292
rect 56953 34588 57069 34616
rect 56953 34532 56983 34588
rect 57039 34532 57069 34588
rect 56953 34508 57069 34532
rect 56953 34452 56983 34508
rect 57039 34452 57069 34508
rect 56953 34428 57069 34452
rect 56953 34372 56983 34428
rect 57039 34372 57069 34428
rect 56953 34348 57069 34372
rect 56953 34292 56983 34348
rect 57039 34292 57069 34348
rect 56953 34264 57069 34292
rect 57795 34588 57911 34616
rect 57795 34532 57825 34588
rect 57881 34532 57911 34588
rect 57795 34508 57911 34532
rect 57795 34452 57825 34508
rect 57881 34452 57911 34508
rect 57795 34428 57911 34452
rect 57795 34372 57825 34428
rect 57881 34372 57911 34428
rect 57795 34348 57911 34372
rect 57795 34292 57825 34348
rect 57881 34292 57911 34348
rect 57795 34264 57911 34292
rect 58461 34588 58525 34616
rect 58461 34532 58465 34588
rect 58521 34532 58525 34588
rect 58461 34508 58525 34532
rect 58461 34452 58465 34508
rect 58521 34452 58525 34508
rect 58461 34428 58525 34452
rect 58461 34372 58465 34428
rect 58521 34372 58525 34428
rect 58461 34348 58525 34372
rect 58461 34292 58465 34348
rect 58521 34292 58525 34348
rect 58461 34264 58525 34292
rect 59018 34588 59134 34616
rect 59018 34532 59048 34588
rect 59104 34532 59134 34588
rect 59018 34508 59134 34532
rect 59018 34452 59048 34508
rect 59104 34452 59134 34508
rect 59018 34428 59134 34452
rect 59018 34372 59048 34428
rect 59104 34372 59134 34428
rect 59018 34348 59134 34372
rect 59018 34292 59048 34348
rect 59104 34292 59134 34348
rect 59018 34264 59134 34292
rect 60296 34588 60412 34616
rect 60296 34532 60326 34588
rect 60382 34532 60412 34588
rect 60296 34508 60412 34532
rect 60296 34452 60326 34508
rect 60382 34452 60412 34508
rect 60296 34428 60412 34452
rect 60296 34372 60326 34428
rect 60382 34372 60412 34428
rect 60296 34348 60412 34372
rect 60296 34292 60326 34348
rect 60382 34292 60412 34348
rect 60296 34264 60412 34292
rect 60454 34588 60570 34616
rect 60454 34532 60484 34588
rect 60540 34532 60570 34588
rect 60454 34508 60570 34532
rect 60454 34452 60484 34508
rect 60540 34452 60570 34508
rect 60454 34428 60570 34452
rect 60454 34372 60484 34428
rect 60540 34372 60570 34428
rect 60454 34348 60570 34372
rect 60454 34292 60484 34348
rect 60540 34292 60570 34348
rect 60454 34264 60570 34292
rect 62509 34588 62683 34616
rect 62509 34532 62528 34588
rect 62584 34532 62608 34588
rect 62664 34532 62683 34588
rect 62509 34508 62683 34532
rect 62509 34452 62528 34508
rect 62584 34452 62608 34508
rect 62664 34452 62683 34508
rect 62509 34428 62683 34452
rect 62509 34372 62528 34428
rect 62584 34372 62608 34428
rect 62664 34372 62683 34428
rect 62509 34348 62683 34372
rect 62509 34292 62528 34348
rect 62584 34292 62608 34348
rect 62664 34292 62683 34348
rect 62509 34264 62683 34292
rect 2152 32236 2352 32264
rect 2152 32180 2184 32236
rect 2240 32180 2264 32236
rect 2320 32180 2352 32236
rect 2152 32156 2352 32180
rect 2152 32100 2184 32156
rect 2240 32100 2264 32156
rect 2320 32100 2352 32156
rect 2152 32076 2352 32100
rect 2152 32020 2184 32076
rect 2240 32020 2264 32076
rect 2320 32020 2352 32076
rect 2152 31996 2352 32020
rect 2152 31940 2184 31996
rect 2240 31940 2264 31996
rect 2320 31940 2352 31996
rect 2152 31912 2352 31940
rect 5374 32236 5468 32264
rect 5374 32180 5393 32236
rect 5449 32180 5468 32236
rect 5374 32156 5468 32180
rect 5374 32100 5393 32156
rect 5449 32100 5468 32156
rect 5374 32076 5468 32100
rect 5374 32020 5393 32076
rect 5449 32020 5468 32076
rect 5374 31996 5468 32020
rect 5374 31940 5393 31996
rect 5449 31940 5468 31996
rect 5374 31912 5468 31940
rect 8264 32236 8358 32264
rect 8264 32180 8283 32236
rect 8339 32180 8358 32236
rect 8264 32156 8358 32180
rect 8264 32100 8283 32156
rect 8339 32100 8358 32156
rect 8264 32076 8358 32100
rect 8264 32020 8283 32076
rect 8339 32020 8358 32076
rect 8264 31996 8358 32020
rect 8264 31940 8283 31996
rect 8339 31940 8358 31996
rect 8264 31912 8358 31940
rect 11154 32236 11248 32264
rect 11154 32180 11173 32236
rect 11229 32180 11248 32236
rect 11154 32156 11248 32180
rect 11154 32100 11173 32156
rect 11229 32100 11248 32156
rect 11154 32076 11248 32100
rect 11154 32020 11173 32076
rect 11229 32020 11248 32076
rect 11154 31996 11248 32020
rect 11154 31940 11173 31996
rect 11229 31940 11248 31996
rect 11154 31912 11248 31940
rect 14044 32236 14138 32264
rect 14044 32180 14063 32236
rect 14119 32180 14138 32236
rect 14044 32156 14138 32180
rect 14044 32100 14063 32156
rect 14119 32100 14138 32156
rect 14044 32076 14138 32100
rect 14044 32020 14063 32076
rect 14119 32020 14138 32076
rect 14044 31996 14138 32020
rect 14044 31940 14063 31996
rect 14119 31940 14138 31996
rect 14044 31912 14138 31940
rect 16934 32236 17028 32264
rect 16934 32180 16953 32236
rect 17009 32180 17028 32236
rect 16934 32156 17028 32180
rect 16934 32100 16953 32156
rect 17009 32100 17028 32156
rect 16934 32076 17028 32100
rect 16934 32020 16953 32076
rect 17009 32020 17028 32076
rect 16934 31996 17028 32020
rect 16934 31940 16953 31996
rect 17009 31940 17028 31996
rect 16934 31912 17028 31940
rect 19824 32236 19918 32264
rect 19824 32180 19843 32236
rect 19899 32180 19918 32236
rect 19824 32156 19918 32180
rect 19824 32100 19843 32156
rect 19899 32100 19918 32156
rect 19824 32076 19918 32100
rect 19824 32020 19843 32076
rect 19899 32020 19918 32076
rect 19824 31996 19918 32020
rect 19824 31940 19843 31996
rect 19899 31940 19918 31996
rect 19824 31912 19918 31940
rect 22714 32236 22808 32264
rect 22714 32180 22733 32236
rect 22789 32180 22808 32236
rect 22714 32156 22808 32180
rect 22714 32100 22733 32156
rect 22789 32100 22808 32156
rect 22714 32076 22808 32100
rect 22714 32020 22733 32076
rect 22789 32020 22808 32076
rect 22714 31996 22808 32020
rect 22714 31940 22733 31996
rect 22789 31940 22808 31996
rect 22714 31912 22808 31940
rect 25604 32236 25698 32264
rect 25604 32180 25623 32236
rect 25679 32180 25698 32236
rect 25604 32156 25698 32180
rect 25604 32100 25623 32156
rect 25679 32100 25698 32156
rect 25604 32076 25698 32100
rect 25604 32020 25623 32076
rect 25679 32020 25698 32076
rect 25604 31996 25698 32020
rect 25604 31940 25623 31996
rect 25679 31940 25698 31996
rect 25604 31912 25698 31940
rect 28494 32236 28588 32264
rect 28494 32180 28513 32236
rect 28569 32180 28588 32236
rect 28494 32156 28588 32180
rect 28494 32100 28513 32156
rect 28569 32100 28588 32156
rect 28494 32076 28588 32100
rect 28494 32020 28513 32076
rect 28569 32020 28588 32076
rect 28494 31996 28588 32020
rect 28494 31940 28513 31996
rect 28569 31940 28588 31996
rect 28494 31912 28588 31940
rect 31384 32236 31478 32264
rect 31384 32180 31403 32236
rect 31459 32180 31478 32236
rect 31384 32156 31478 32180
rect 31384 32100 31403 32156
rect 31459 32100 31478 32156
rect 31384 32076 31478 32100
rect 31384 32020 31403 32076
rect 31459 32020 31478 32076
rect 31384 31996 31478 32020
rect 31384 31940 31403 31996
rect 31459 31940 31478 31996
rect 31384 31912 31478 31940
rect 34274 32236 34368 32264
rect 34274 32180 34293 32236
rect 34349 32180 34368 32236
rect 34274 32156 34368 32180
rect 34274 32100 34293 32156
rect 34349 32100 34368 32156
rect 34274 32076 34368 32100
rect 34274 32020 34293 32076
rect 34349 32020 34368 32076
rect 34274 31996 34368 32020
rect 34274 31940 34293 31996
rect 34349 31940 34368 31996
rect 34274 31912 34368 31940
rect 37164 32236 37258 32264
rect 37164 32180 37183 32236
rect 37239 32180 37258 32236
rect 37164 32156 37258 32180
rect 37164 32100 37183 32156
rect 37239 32100 37258 32156
rect 37164 32076 37258 32100
rect 37164 32020 37183 32076
rect 37239 32020 37258 32076
rect 37164 31996 37258 32020
rect 37164 31940 37183 31996
rect 37239 31940 37258 31996
rect 37164 31912 37258 31940
rect 40054 32236 40148 32264
rect 40054 32180 40073 32236
rect 40129 32180 40148 32236
rect 40054 32156 40148 32180
rect 40054 32100 40073 32156
rect 40129 32100 40148 32156
rect 40054 32076 40148 32100
rect 40054 32020 40073 32076
rect 40129 32020 40148 32076
rect 40054 31996 40148 32020
rect 40054 31940 40073 31996
rect 40129 31940 40148 31996
rect 40054 31912 40148 31940
rect 42944 32236 43038 32264
rect 42944 32180 42963 32236
rect 43019 32180 43038 32236
rect 42944 32156 43038 32180
rect 42944 32100 42963 32156
rect 43019 32100 43038 32156
rect 42944 32076 43038 32100
rect 42944 32020 42963 32076
rect 43019 32020 43038 32076
rect 42944 31996 43038 32020
rect 42944 31940 42963 31996
rect 43019 31940 43038 31996
rect 42944 31912 43038 31940
rect 45834 32236 45928 32264
rect 45834 32180 45853 32236
rect 45909 32180 45928 32236
rect 45834 32156 45928 32180
rect 45834 32100 45853 32156
rect 45909 32100 45928 32156
rect 45834 32076 45928 32100
rect 45834 32020 45853 32076
rect 45909 32020 45928 32076
rect 45834 31996 45928 32020
rect 45834 31940 45853 31996
rect 45909 31940 45928 31996
rect 45834 31912 45928 31940
rect 48781 32236 48875 32264
rect 48781 32180 48800 32236
rect 48856 32180 48875 32236
rect 48781 32156 48875 32180
rect 48781 32100 48800 32156
rect 48856 32100 48875 32156
rect 48781 32076 48875 32100
rect 48781 32020 48800 32076
rect 48856 32020 48875 32076
rect 48781 31996 48875 32020
rect 48781 31940 48800 31996
rect 48856 31940 48875 31996
rect 48781 31912 48875 31940
rect 49630 32236 49830 32264
rect 49630 32180 49662 32236
rect 49718 32180 49742 32236
rect 49798 32180 49830 32236
rect 49630 32156 49830 32180
rect 49630 32100 49662 32156
rect 49718 32100 49742 32156
rect 49798 32100 49830 32156
rect 49630 32076 49830 32100
rect 49630 32020 49662 32076
rect 49718 32020 49742 32076
rect 49798 32020 49830 32076
rect 49630 31996 49830 32020
rect 49630 31940 49662 31996
rect 49718 31940 49742 31996
rect 49798 31940 49830 31996
rect 49630 31912 49830 31940
rect 52920 32236 53048 32264
rect 52920 32180 52956 32236
rect 53012 32180 53048 32236
rect 52920 32156 53048 32180
rect 52920 32100 52956 32156
rect 53012 32100 53048 32156
rect 52920 32076 53048 32100
rect 52920 32020 52956 32076
rect 53012 32020 53048 32076
rect 52920 31996 53048 32020
rect 52920 31940 52956 31996
rect 53012 31940 53048 31996
rect 52920 31912 53048 31940
rect 53078 32236 53206 32264
rect 53078 32180 53114 32236
rect 53170 32180 53206 32236
rect 53078 32156 53206 32180
rect 53078 32100 53114 32156
rect 53170 32100 53206 32156
rect 53078 32076 53206 32100
rect 53078 32020 53114 32076
rect 53170 32020 53206 32076
rect 53078 31996 53206 32020
rect 53078 31940 53114 31996
rect 53170 31940 53206 31996
rect 53078 31912 53206 31940
rect 53434 32236 53562 32264
rect 53434 32180 53470 32236
rect 53526 32180 53562 32236
rect 53434 32156 53562 32180
rect 53434 32100 53470 32156
rect 53526 32100 53562 32156
rect 53434 32076 53562 32100
rect 53434 32020 53470 32076
rect 53526 32020 53562 32076
rect 53434 31996 53562 32020
rect 53434 31940 53470 31996
rect 53526 31940 53562 31996
rect 53434 31912 53562 31940
rect 54752 32236 54880 32264
rect 54752 32180 54788 32236
rect 54844 32180 54880 32236
rect 54752 32156 54880 32180
rect 54752 32100 54788 32156
rect 54844 32100 54880 32156
rect 54752 32076 54880 32100
rect 54752 32020 54788 32076
rect 54844 32020 54880 32076
rect 54752 31996 54880 32020
rect 54752 31940 54788 31996
rect 54844 31940 54880 31996
rect 54752 31912 54880 31940
rect 55345 32236 55473 32264
rect 55345 32180 55381 32236
rect 55437 32180 55473 32236
rect 55345 32156 55473 32180
rect 55345 32100 55381 32156
rect 55437 32100 55473 32156
rect 55345 32076 55473 32100
rect 55345 32020 55381 32076
rect 55437 32020 55473 32076
rect 55345 31996 55473 32020
rect 55345 31940 55381 31996
rect 55437 31940 55473 31996
rect 55345 31912 55473 31940
rect 56491 32236 56619 32264
rect 56491 32180 56527 32236
rect 56583 32180 56619 32236
rect 56491 32156 56619 32180
rect 56491 32100 56527 32156
rect 56583 32100 56619 32156
rect 56491 32076 56619 32100
rect 56491 32020 56527 32076
rect 56583 32020 56619 32076
rect 56491 31996 56619 32020
rect 56491 31940 56527 31996
rect 56583 31940 56619 31996
rect 56491 31912 56619 31940
rect 57941 32236 58121 32264
rect 57941 32180 57963 32236
rect 58019 32180 58043 32236
rect 58099 32180 58121 32236
rect 57941 32156 58121 32180
rect 57941 32100 57963 32156
rect 58019 32100 58043 32156
rect 58099 32100 58121 32156
rect 57941 32076 58121 32100
rect 57941 32020 57963 32076
rect 58019 32020 58043 32076
rect 58099 32020 58121 32076
rect 57941 31996 58121 32020
rect 57941 31940 57963 31996
rect 58019 31940 58043 31996
rect 58099 31940 58121 31996
rect 57941 31912 58121 31940
rect 59164 32236 59304 32264
rect 59164 32180 59206 32236
rect 59262 32180 59304 32236
rect 59164 32156 59304 32180
rect 59164 32100 59206 32156
rect 59262 32100 59304 32156
rect 59164 32076 59304 32100
rect 59164 32020 59206 32076
rect 59262 32020 59304 32076
rect 59164 31996 59304 32020
rect 59164 31940 59206 31996
rect 59262 31940 59304 31996
rect 59164 31912 59304 31940
rect 59334 32236 59450 32264
rect 59334 32180 59364 32236
rect 59420 32180 59450 32236
rect 59334 32156 59450 32180
rect 59334 32100 59364 32156
rect 59420 32100 59450 32156
rect 59334 32076 59450 32100
rect 59334 32020 59364 32076
rect 59420 32020 59450 32076
rect 59334 31996 59450 32020
rect 59334 31940 59364 31996
rect 59420 31940 59450 31996
rect 59334 31912 59450 31940
rect 59642 32236 59758 32264
rect 59642 32180 59672 32236
rect 59728 32180 59758 32236
rect 59642 32156 59758 32180
rect 59642 32100 59672 32156
rect 59728 32100 59758 32156
rect 59642 32076 59758 32100
rect 59642 32020 59672 32076
rect 59728 32020 59758 32076
rect 59642 31996 59758 32020
rect 59642 31940 59672 31996
rect 59728 31940 59758 31996
rect 59642 31912 59758 31940
rect 59788 32236 59904 32264
rect 59788 32180 59818 32236
rect 59874 32180 59904 32236
rect 59788 32156 59904 32180
rect 59788 32100 59818 32156
rect 59874 32100 59904 32156
rect 59788 32076 59904 32100
rect 59788 32020 59818 32076
rect 59874 32020 59904 32076
rect 59788 31996 59904 32020
rect 59788 31940 59818 31996
rect 59874 31940 59904 31996
rect 59788 31912 59904 31940
rect 59934 32236 60110 32264
rect 59934 32180 59954 32236
rect 60010 32180 60034 32236
rect 60090 32180 60110 32236
rect 59934 32156 60110 32180
rect 59934 32100 59954 32156
rect 60010 32100 60034 32156
rect 60090 32100 60110 32156
rect 59934 32076 60110 32100
rect 59934 32020 59954 32076
rect 60010 32020 60034 32076
rect 60090 32020 60110 32076
rect 59934 31996 60110 32020
rect 59934 31940 59954 31996
rect 60010 31940 60034 31996
rect 60090 31940 60110 31996
rect 59934 31912 60110 31940
rect 62307 32236 62481 32264
rect 62307 32180 62326 32236
rect 62382 32180 62406 32236
rect 62462 32180 62481 32236
rect 62307 32156 62481 32180
rect 62307 32100 62326 32156
rect 62382 32100 62406 32156
rect 62462 32100 62481 32156
rect 62307 32076 62481 32100
rect 62307 32020 62326 32076
rect 62382 32020 62406 32076
rect 62462 32020 62481 32076
rect 62307 31996 62481 32020
rect 62307 31940 62326 31996
rect 62382 31940 62406 31996
rect 62462 31940 62481 31996
rect 62307 31912 62481 31940
rect 2020 24588 2124 24616
rect 2020 24532 2044 24588
rect 2100 24532 2124 24588
rect 2020 24508 2124 24532
rect 2020 24452 2044 24508
rect 2100 24452 2124 24508
rect 2020 24428 2124 24452
rect 2020 24372 2044 24428
rect 2100 24372 2124 24428
rect 2020 24348 2124 24372
rect 2020 24292 2044 24348
rect 2100 24292 2124 24348
rect 2020 24264 2124 24292
rect 5521 24588 5615 24616
rect 5521 24532 5540 24588
rect 5596 24532 5615 24588
rect 5521 24508 5615 24532
rect 5521 24452 5540 24508
rect 5596 24452 5615 24508
rect 5521 24428 5615 24452
rect 5521 24372 5540 24428
rect 5596 24372 5615 24428
rect 5521 24348 5615 24372
rect 5521 24292 5540 24348
rect 5596 24292 5615 24348
rect 5521 24264 5615 24292
rect 8411 24588 8505 24616
rect 8411 24532 8430 24588
rect 8486 24532 8505 24588
rect 8411 24508 8505 24532
rect 8411 24452 8430 24508
rect 8486 24452 8505 24508
rect 8411 24428 8505 24452
rect 8411 24372 8430 24428
rect 8486 24372 8505 24428
rect 8411 24348 8505 24372
rect 8411 24292 8430 24348
rect 8486 24292 8505 24348
rect 8411 24264 8505 24292
rect 11301 24588 11395 24616
rect 11301 24532 11320 24588
rect 11376 24532 11395 24588
rect 11301 24508 11395 24532
rect 11301 24452 11320 24508
rect 11376 24452 11395 24508
rect 11301 24428 11395 24452
rect 11301 24372 11320 24428
rect 11376 24372 11395 24428
rect 11301 24348 11395 24372
rect 11301 24292 11320 24348
rect 11376 24292 11395 24348
rect 11301 24264 11395 24292
rect 14191 24588 14285 24616
rect 14191 24532 14210 24588
rect 14266 24532 14285 24588
rect 14191 24508 14285 24532
rect 14191 24452 14210 24508
rect 14266 24452 14285 24508
rect 14191 24428 14285 24452
rect 14191 24372 14210 24428
rect 14266 24372 14285 24428
rect 14191 24348 14285 24372
rect 14191 24292 14210 24348
rect 14266 24292 14285 24348
rect 14191 24264 14285 24292
rect 17081 24588 17175 24616
rect 17081 24532 17100 24588
rect 17156 24532 17175 24588
rect 17081 24508 17175 24532
rect 17081 24452 17100 24508
rect 17156 24452 17175 24508
rect 17081 24428 17175 24452
rect 17081 24372 17100 24428
rect 17156 24372 17175 24428
rect 17081 24348 17175 24372
rect 17081 24292 17100 24348
rect 17156 24292 17175 24348
rect 17081 24264 17175 24292
rect 19971 24588 20065 24616
rect 19971 24532 19990 24588
rect 20046 24532 20065 24588
rect 19971 24508 20065 24532
rect 19971 24452 19990 24508
rect 20046 24452 20065 24508
rect 19971 24428 20065 24452
rect 19971 24372 19990 24428
rect 20046 24372 20065 24428
rect 19971 24348 20065 24372
rect 19971 24292 19990 24348
rect 20046 24292 20065 24348
rect 19971 24264 20065 24292
rect 22861 24588 22955 24616
rect 22861 24532 22880 24588
rect 22936 24532 22955 24588
rect 22861 24508 22955 24532
rect 22861 24452 22880 24508
rect 22936 24452 22955 24508
rect 22861 24428 22955 24452
rect 22861 24372 22880 24428
rect 22936 24372 22955 24428
rect 22861 24348 22955 24372
rect 22861 24292 22880 24348
rect 22936 24292 22955 24348
rect 22861 24264 22955 24292
rect 25751 24588 25845 24616
rect 25751 24532 25770 24588
rect 25826 24532 25845 24588
rect 25751 24508 25845 24532
rect 25751 24452 25770 24508
rect 25826 24452 25845 24508
rect 25751 24428 25845 24452
rect 25751 24372 25770 24428
rect 25826 24372 25845 24428
rect 25751 24348 25845 24372
rect 25751 24292 25770 24348
rect 25826 24292 25845 24348
rect 25751 24264 25845 24292
rect 28641 24588 28735 24616
rect 28641 24532 28660 24588
rect 28716 24532 28735 24588
rect 28641 24508 28735 24532
rect 28641 24452 28660 24508
rect 28716 24452 28735 24508
rect 28641 24428 28735 24452
rect 28641 24372 28660 24428
rect 28716 24372 28735 24428
rect 28641 24348 28735 24372
rect 28641 24292 28660 24348
rect 28716 24292 28735 24348
rect 28641 24264 28735 24292
rect 31531 24588 31625 24616
rect 31531 24532 31550 24588
rect 31606 24532 31625 24588
rect 31531 24508 31625 24532
rect 31531 24452 31550 24508
rect 31606 24452 31625 24508
rect 31531 24428 31625 24452
rect 31531 24372 31550 24428
rect 31606 24372 31625 24428
rect 31531 24348 31625 24372
rect 31531 24292 31550 24348
rect 31606 24292 31625 24348
rect 31531 24264 31625 24292
rect 34421 24588 34515 24616
rect 34421 24532 34440 24588
rect 34496 24532 34515 24588
rect 34421 24508 34515 24532
rect 34421 24452 34440 24508
rect 34496 24452 34515 24508
rect 34421 24428 34515 24452
rect 34421 24372 34440 24428
rect 34496 24372 34515 24428
rect 34421 24348 34515 24372
rect 34421 24292 34440 24348
rect 34496 24292 34515 24348
rect 34421 24264 34515 24292
rect 37311 24588 37405 24616
rect 37311 24532 37330 24588
rect 37386 24532 37405 24588
rect 37311 24508 37405 24532
rect 37311 24452 37330 24508
rect 37386 24452 37405 24508
rect 37311 24428 37405 24452
rect 37311 24372 37330 24428
rect 37386 24372 37405 24428
rect 37311 24348 37405 24372
rect 37311 24292 37330 24348
rect 37386 24292 37405 24348
rect 37311 24264 37405 24292
rect 40201 24588 40295 24616
rect 40201 24532 40220 24588
rect 40276 24532 40295 24588
rect 40201 24508 40295 24532
rect 40201 24452 40220 24508
rect 40276 24452 40295 24508
rect 40201 24428 40295 24452
rect 40201 24372 40220 24428
rect 40276 24372 40295 24428
rect 40201 24348 40295 24372
rect 40201 24292 40220 24348
rect 40276 24292 40295 24348
rect 40201 24264 40295 24292
rect 43091 24588 43185 24616
rect 43091 24532 43110 24588
rect 43166 24532 43185 24588
rect 43091 24508 43185 24532
rect 43091 24452 43110 24508
rect 43166 24452 43185 24508
rect 43091 24428 43185 24452
rect 43091 24372 43110 24428
rect 43166 24372 43185 24428
rect 43091 24348 43185 24372
rect 43091 24292 43110 24348
rect 43166 24292 43185 24348
rect 43091 24264 43185 24292
rect 45981 24588 46075 24616
rect 45981 24532 46000 24588
rect 46056 24532 46075 24588
rect 45981 24508 46075 24532
rect 45981 24452 46000 24508
rect 46056 24452 46075 24508
rect 45981 24428 46075 24452
rect 45981 24372 46000 24428
rect 46056 24372 46075 24428
rect 45981 24348 46075 24372
rect 45981 24292 46000 24348
rect 46056 24292 46075 24348
rect 45981 24264 46075 24292
rect 48989 24588 49083 24616
rect 48989 24532 49008 24588
rect 49064 24532 49083 24588
rect 48989 24508 49083 24532
rect 48989 24452 49008 24508
rect 49064 24452 49083 24508
rect 48989 24428 49083 24452
rect 48989 24372 49008 24428
rect 49064 24372 49083 24428
rect 48989 24348 49083 24372
rect 48989 24292 49008 24348
rect 49064 24292 49083 24348
rect 48989 24264 49083 24292
rect 52210 24588 52320 24616
rect 52210 24532 52237 24588
rect 52293 24532 52320 24588
rect 52210 24508 52320 24532
rect 52210 24452 52237 24508
rect 52293 24452 52320 24508
rect 52210 24428 52320 24452
rect 52210 24372 52237 24428
rect 52293 24372 52320 24428
rect 52210 24348 52320 24372
rect 52210 24292 52237 24348
rect 52293 24292 52320 24348
rect 52210 24264 52320 24292
rect 53602 24588 53730 24616
rect 53602 24532 53638 24588
rect 53694 24532 53730 24588
rect 53602 24508 53730 24532
rect 53602 24452 53638 24508
rect 53694 24452 53730 24508
rect 53602 24428 53730 24452
rect 53602 24372 53638 24428
rect 53694 24372 53730 24428
rect 53602 24348 53730 24372
rect 53602 24292 53638 24348
rect 53694 24292 53730 24348
rect 53602 24264 53730 24292
rect 53770 24588 53898 24616
rect 53770 24532 53806 24588
rect 53862 24532 53898 24588
rect 53770 24508 53898 24532
rect 53770 24452 53806 24508
rect 53862 24452 53898 24508
rect 53770 24428 53898 24452
rect 53770 24372 53806 24428
rect 53862 24372 53898 24428
rect 53770 24348 53898 24372
rect 53770 24292 53806 24348
rect 53862 24292 53898 24348
rect 53770 24264 53898 24292
rect 54514 24588 54642 24616
rect 54514 24532 54550 24588
rect 54606 24532 54642 24588
rect 54514 24508 54642 24532
rect 54514 24452 54550 24508
rect 54606 24452 54642 24508
rect 54514 24428 54642 24452
rect 54514 24372 54550 24428
rect 54606 24372 54642 24428
rect 54514 24348 54642 24372
rect 54514 24292 54550 24348
rect 54606 24292 54642 24348
rect 54514 24264 54642 24292
rect 54910 24588 55026 24616
rect 54910 24532 54940 24588
rect 54996 24532 55026 24588
rect 54910 24508 55026 24532
rect 54910 24452 54940 24508
rect 54996 24452 55026 24508
rect 54910 24428 55026 24452
rect 54910 24372 54940 24428
rect 54996 24372 55026 24428
rect 54910 24348 55026 24372
rect 54910 24292 54940 24348
rect 54996 24292 55026 24348
rect 54910 24264 55026 24292
rect 55620 24588 55748 24616
rect 55620 24532 55656 24588
rect 55712 24532 55748 24588
rect 55620 24508 55748 24532
rect 55620 24452 55656 24508
rect 55712 24452 55748 24508
rect 55620 24428 55748 24452
rect 55620 24372 55656 24428
rect 55712 24372 55748 24428
rect 55620 24348 55748 24372
rect 55620 24292 55656 24348
rect 55712 24292 55748 24348
rect 55620 24264 55748 24292
rect 56198 24588 56326 24616
rect 56198 24532 56234 24588
rect 56290 24532 56326 24588
rect 56198 24508 56326 24532
rect 56198 24452 56234 24508
rect 56290 24452 56326 24508
rect 56198 24428 56326 24452
rect 56198 24372 56234 24428
rect 56290 24372 56326 24428
rect 56198 24348 56326 24372
rect 56198 24292 56234 24348
rect 56290 24292 56326 24348
rect 56198 24264 56326 24292
rect 56649 24588 56765 24616
rect 56649 24532 56679 24588
rect 56735 24532 56765 24588
rect 56649 24508 56765 24532
rect 56649 24452 56679 24508
rect 56735 24452 56765 24508
rect 56649 24428 56765 24452
rect 56649 24372 56679 24428
rect 56735 24372 56765 24428
rect 56649 24348 56765 24372
rect 56649 24292 56679 24348
rect 56735 24292 56765 24348
rect 56649 24264 56765 24292
rect 56953 24588 57069 24616
rect 56953 24532 56983 24588
rect 57039 24532 57069 24588
rect 56953 24508 57069 24532
rect 56953 24452 56983 24508
rect 57039 24452 57069 24508
rect 56953 24428 57069 24452
rect 56953 24372 56983 24428
rect 57039 24372 57069 24428
rect 56953 24348 57069 24372
rect 56953 24292 56983 24348
rect 57039 24292 57069 24348
rect 56953 24264 57069 24292
rect 57795 24588 57911 24616
rect 57795 24532 57825 24588
rect 57881 24532 57911 24588
rect 57795 24508 57911 24532
rect 57795 24452 57825 24508
rect 57881 24452 57911 24508
rect 57795 24428 57911 24452
rect 57795 24372 57825 24428
rect 57881 24372 57911 24428
rect 57795 24348 57911 24372
rect 57795 24292 57825 24348
rect 57881 24292 57911 24348
rect 57795 24264 57911 24292
rect 58461 24588 58525 24616
rect 58461 24532 58465 24588
rect 58521 24532 58525 24588
rect 58461 24508 58525 24532
rect 58461 24452 58465 24508
rect 58521 24452 58525 24508
rect 58461 24428 58525 24452
rect 58461 24372 58465 24428
rect 58521 24372 58525 24428
rect 58461 24348 58525 24372
rect 58461 24292 58465 24348
rect 58521 24292 58525 24348
rect 58461 24264 58525 24292
rect 59018 24588 59134 24616
rect 59018 24532 59048 24588
rect 59104 24532 59134 24588
rect 59018 24508 59134 24532
rect 59018 24452 59048 24508
rect 59104 24452 59134 24508
rect 59018 24428 59134 24452
rect 59018 24372 59048 24428
rect 59104 24372 59134 24428
rect 59018 24348 59134 24372
rect 59018 24292 59048 24348
rect 59104 24292 59134 24348
rect 59018 24264 59134 24292
rect 60296 24588 60412 24616
rect 60296 24532 60326 24588
rect 60382 24532 60412 24588
rect 60296 24508 60412 24532
rect 60296 24452 60326 24508
rect 60382 24452 60412 24508
rect 60296 24428 60412 24452
rect 60296 24372 60326 24428
rect 60382 24372 60412 24428
rect 60296 24348 60412 24372
rect 60296 24292 60326 24348
rect 60382 24292 60412 24348
rect 60296 24264 60412 24292
rect 60454 24588 60570 24616
rect 60454 24532 60484 24588
rect 60540 24532 60570 24588
rect 60454 24508 60570 24532
rect 60454 24452 60484 24508
rect 60540 24452 60570 24508
rect 60454 24428 60570 24452
rect 60454 24372 60484 24428
rect 60540 24372 60570 24428
rect 60454 24348 60570 24372
rect 60454 24292 60484 24348
rect 60540 24292 60570 24348
rect 60454 24264 60570 24292
rect 62509 24588 62683 24616
rect 62509 24532 62528 24588
rect 62584 24532 62608 24588
rect 62664 24532 62683 24588
rect 62509 24508 62683 24532
rect 62509 24452 62528 24508
rect 62584 24452 62608 24508
rect 62664 24452 62683 24508
rect 62509 24428 62683 24452
rect 62509 24372 62528 24428
rect 62584 24372 62608 24428
rect 62664 24372 62683 24428
rect 62509 24348 62683 24372
rect 62509 24292 62528 24348
rect 62584 24292 62608 24348
rect 62664 24292 62683 24348
rect 62509 24264 62683 24292
rect 2152 22236 2352 22264
rect 2152 22180 2184 22236
rect 2240 22180 2264 22236
rect 2320 22180 2352 22236
rect 2152 22156 2352 22180
rect 2152 22100 2184 22156
rect 2240 22100 2264 22156
rect 2320 22100 2352 22156
rect 2152 22076 2352 22100
rect 2152 22020 2184 22076
rect 2240 22020 2264 22076
rect 2320 22020 2352 22076
rect 2152 21996 2352 22020
rect 2152 21940 2184 21996
rect 2240 21940 2264 21996
rect 2320 21940 2352 21996
rect 2152 21912 2352 21940
rect 5374 22236 5468 22264
rect 5374 22180 5393 22236
rect 5449 22180 5468 22236
rect 5374 22156 5468 22180
rect 5374 22100 5393 22156
rect 5449 22100 5468 22156
rect 5374 22076 5468 22100
rect 5374 22020 5393 22076
rect 5449 22020 5468 22076
rect 5374 21996 5468 22020
rect 5374 21940 5393 21996
rect 5449 21940 5468 21996
rect 5374 21912 5468 21940
rect 8264 22236 8358 22264
rect 8264 22180 8283 22236
rect 8339 22180 8358 22236
rect 8264 22156 8358 22180
rect 8264 22100 8283 22156
rect 8339 22100 8358 22156
rect 8264 22076 8358 22100
rect 8264 22020 8283 22076
rect 8339 22020 8358 22076
rect 8264 21996 8358 22020
rect 8264 21940 8283 21996
rect 8339 21940 8358 21996
rect 8264 21912 8358 21940
rect 11154 22236 11248 22264
rect 11154 22180 11173 22236
rect 11229 22180 11248 22236
rect 11154 22156 11248 22180
rect 11154 22100 11173 22156
rect 11229 22100 11248 22156
rect 11154 22076 11248 22100
rect 11154 22020 11173 22076
rect 11229 22020 11248 22076
rect 11154 21996 11248 22020
rect 11154 21940 11173 21996
rect 11229 21940 11248 21996
rect 11154 21912 11248 21940
rect 14044 22236 14138 22264
rect 14044 22180 14063 22236
rect 14119 22180 14138 22236
rect 14044 22156 14138 22180
rect 14044 22100 14063 22156
rect 14119 22100 14138 22156
rect 14044 22076 14138 22100
rect 14044 22020 14063 22076
rect 14119 22020 14138 22076
rect 14044 21996 14138 22020
rect 14044 21940 14063 21996
rect 14119 21940 14138 21996
rect 14044 21912 14138 21940
rect 16934 22236 17028 22264
rect 16934 22180 16953 22236
rect 17009 22180 17028 22236
rect 16934 22156 17028 22180
rect 16934 22100 16953 22156
rect 17009 22100 17028 22156
rect 16934 22076 17028 22100
rect 16934 22020 16953 22076
rect 17009 22020 17028 22076
rect 16934 21996 17028 22020
rect 16934 21940 16953 21996
rect 17009 21940 17028 21996
rect 16934 21912 17028 21940
rect 19824 22236 19918 22264
rect 19824 22180 19843 22236
rect 19899 22180 19918 22236
rect 19824 22156 19918 22180
rect 19824 22100 19843 22156
rect 19899 22100 19918 22156
rect 19824 22076 19918 22100
rect 19824 22020 19843 22076
rect 19899 22020 19918 22076
rect 19824 21996 19918 22020
rect 19824 21940 19843 21996
rect 19899 21940 19918 21996
rect 19824 21912 19918 21940
rect 22714 22236 22808 22264
rect 22714 22180 22733 22236
rect 22789 22180 22808 22236
rect 22714 22156 22808 22180
rect 22714 22100 22733 22156
rect 22789 22100 22808 22156
rect 22714 22076 22808 22100
rect 22714 22020 22733 22076
rect 22789 22020 22808 22076
rect 22714 21996 22808 22020
rect 22714 21940 22733 21996
rect 22789 21940 22808 21996
rect 22714 21912 22808 21940
rect 25604 22236 25698 22264
rect 25604 22180 25623 22236
rect 25679 22180 25698 22236
rect 25604 22156 25698 22180
rect 25604 22100 25623 22156
rect 25679 22100 25698 22156
rect 25604 22076 25698 22100
rect 25604 22020 25623 22076
rect 25679 22020 25698 22076
rect 25604 21996 25698 22020
rect 25604 21940 25623 21996
rect 25679 21940 25698 21996
rect 25604 21912 25698 21940
rect 28494 22236 28588 22264
rect 28494 22180 28513 22236
rect 28569 22180 28588 22236
rect 28494 22156 28588 22180
rect 28494 22100 28513 22156
rect 28569 22100 28588 22156
rect 28494 22076 28588 22100
rect 28494 22020 28513 22076
rect 28569 22020 28588 22076
rect 28494 21996 28588 22020
rect 28494 21940 28513 21996
rect 28569 21940 28588 21996
rect 28494 21912 28588 21940
rect 31384 22236 31478 22264
rect 31384 22180 31403 22236
rect 31459 22180 31478 22236
rect 31384 22156 31478 22180
rect 31384 22100 31403 22156
rect 31459 22100 31478 22156
rect 31384 22076 31478 22100
rect 31384 22020 31403 22076
rect 31459 22020 31478 22076
rect 31384 21996 31478 22020
rect 31384 21940 31403 21996
rect 31459 21940 31478 21996
rect 31384 21912 31478 21940
rect 34274 22236 34368 22264
rect 34274 22180 34293 22236
rect 34349 22180 34368 22236
rect 34274 22156 34368 22180
rect 34274 22100 34293 22156
rect 34349 22100 34368 22156
rect 34274 22076 34368 22100
rect 34274 22020 34293 22076
rect 34349 22020 34368 22076
rect 34274 21996 34368 22020
rect 34274 21940 34293 21996
rect 34349 21940 34368 21996
rect 34274 21912 34368 21940
rect 37164 22236 37258 22264
rect 37164 22180 37183 22236
rect 37239 22180 37258 22236
rect 37164 22156 37258 22180
rect 37164 22100 37183 22156
rect 37239 22100 37258 22156
rect 37164 22076 37258 22100
rect 37164 22020 37183 22076
rect 37239 22020 37258 22076
rect 37164 21996 37258 22020
rect 37164 21940 37183 21996
rect 37239 21940 37258 21996
rect 37164 21912 37258 21940
rect 40054 22236 40148 22264
rect 40054 22180 40073 22236
rect 40129 22180 40148 22236
rect 40054 22156 40148 22180
rect 40054 22100 40073 22156
rect 40129 22100 40148 22156
rect 40054 22076 40148 22100
rect 40054 22020 40073 22076
rect 40129 22020 40148 22076
rect 40054 21996 40148 22020
rect 40054 21940 40073 21996
rect 40129 21940 40148 21996
rect 40054 21912 40148 21940
rect 42944 22236 43038 22264
rect 42944 22180 42963 22236
rect 43019 22180 43038 22236
rect 42944 22156 43038 22180
rect 42944 22100 42963 22156
rect 43019 22100 43038 22156
rect 42944 22076 43038 22100
rect 42944 22020 42963 22076
rect 43019 22020 43038 22076
rect 42944 21996 43038 22020
rect 42944 21940 42963 21996
rect 43019 21940 43038 21996
rect 42944 21912 43038 21940
rect 45834 22236 45928 22264
rect 45834 22180 45853 22236
rect 45909 22180 45928 22236
rect 45834 22156 45928 22180
rect 45834 22100 45853 22156
rect 45909 22100 45928 22156
rect 45834 22076 45928 22100
rect 45834 22020 45853 22076
rect 45909 22020 45928 22076
rect 45834 21996 45928 22020
rect 45834 21940 45853 21996
rect 45909 21940 45928 21996
rect 45834 21912 45928 21940
rect 48781 22236 48875 22264
rect 48781 22180 48800 22236
rect 48856 22180 48875 22236
rect 48781 22156 48875 22180
rect 48781 22100 48800 22156
rect 48856 22100 48875 22156
rect 48781 22076 48875 22100
rect 48781 22020 48800 22076
rect 48856 22020 48875 22076
rect 48781 21996 48875 22020
rect 48781 21940 48800 21996
rect 48856 21940 48875 21996
rect 48781 21912 48875 21940
rect 49630 22236 49830 22264
rect 49630 22180 49662 22236
rect 49718 22180 49742 22236
rect 49798 22180 49830 22236
rect 49630 22156 49830 22180
rect 49630 22100 49662 22156
rect 49718 22100 49742 22156
rect 49798 22100 49830 22156
rect 49630 22076 49830 22100
rect 49630 22020 49662 22076
rect 49718 22020 49742 22076
rect 49798 22020 49830 22076
rect 49630 21996 49830 22020
rect 49630 21940 49662 21996
rect 49718 21940 49742 21996
rect 49798 21940 49830 21996
rect 49630 21912 49830 21940
rect 52920 22236 53048 22264
rect 52920 22180 52956 22236
rect 53012 22180 53048 22236
rect 52920 22156 53048 22180
rect 52920 22100 52956 22156
rect 53012 22100 53048 22156
rect 52920 22076 53048 22100
rect 52920 22020 52956 22076
rect 53012 22020 53048 22076
rect 52920 21996 53048 22020
rect 52920 21940 52956 21996
rect 53012 21940 53048 21996
rect 52920 21912 53048 21940
rect 53078 22236 53206 22264
rect 53078 22180 53114 22236
rect 53170 22180 53206 22236
rect 53078 22156 53206 22180
rect 53078 22100 53114 22156
rect 53170 22100 53206 22156
rect 53078 22076 53206 22100
rect 53078 22020 53114 22076
rect 53170 22020 53206 22076
rect 53078 21996 53206 22020
rect 53078 21940 53114 21996
rect 53170 21940 53206 21996
rect 53078 21912 53206 21940
rect 53434 22236 53562 22264
rect 53434 22180 53470 22236
rect 53526 22180 53562 22236
rect 53434 22156 53562 22180
rect 53434 22100 53470 22156
rect 53526 22100 53562 22156
rect 53434 22076 53562 22100
rect 53434 22020 53470 22076
rect 53526 22020 53562 22076
rect 53434 21996 53562 22020
rect 53434 21940 53470 21996
rect 53526 21940 53562 21996
rect 53434 21912 53562 21940
rect 54752 22236 54880 22264
rect 54752 22180 54788 22236
rect 54844 22180 54880 22236
rect 54752 22156 54880 22180
rect 54752 22100 54788 22156
rect 54844 22100 54880 22156
rect 54752 22076 54880 22100
rect 54752 22020 54788 22076
rect 54844 22020 54880 22076
rect 54752 21996 54880 22020
rect 54752 21940 54788 21996
rect 54844 21940 54880 21996
rect 54752 21912 54880 21940
rect 55345 22236 55473 22264
rect 55345 22180 55381 22236
rect 55437 22180 55473 22236
rect 55345 22156 55473 22180
rect 55345 22100 55381 22156
rect 55437 22100 55473 22156
rect 55345 22076 55473 22100
rect 55345 22020 55381 22076
rect 55437 22020 55473 22076
rect 55345 21996 55473 22020
rect 55345 21940 55381 21996
rect 55437 21940 55473 21996
rect 55345 21912 55473 21940
rect 56491 22236 56619 22264
rect 56491 22180 56527 22236
rect 56583 22180 56619 22236
rect 56491 22156 56619 22180
rect 56491 22100 56527 22156
rect 56583 22100 56619 22156
rect 56491 22076 56619 22100
rect 56491 22020 56527 22076
rect 56583 22020 56619 22076
rect 56491 21996 56619 22020
rect 56491 21940 56527 21996
rect 56583 21940 56619 21996
rect 56491 21912 56619 21940
rect 57941 22236 58121 22264
rect 57941 22180 57963 22236
rect 58019 22180 58043 22236
rect 58099 22180 58121 22236
rect 57941 22156 58121 22180
rect 57941 22100 57963 22156
rect 58019 22100 58043 22156
rect 58099 22100 58121 22156
rect 57941 22076 58121 22100
rect 57941 22020 57963 22076
rect 58019 22020 58043 22076
rect 58099 22020 58121 22076
rect 57941 21996 58121 22020
rect 57941 21940 57963 21996
rect 58019 21940 58043 21996
rect 58099 21940 58121 21996
rect 57941 21912 58121 21940
rect 59164 22236 59304 22264
rect 59164 22180 59206 22236
rect 59262 22180 59304 22236
rect 59164 22156 59304 22180
rect 59164 22100 59206 22156
rect 59262 22100 59304 22156
rect 59164 22076 59304 22100
rect 59164 22020 59206 22076
rect 59262 22020 59304 22076
rect 59164 21996 59304 22020
rect 59164 21940 59206 21996
rect 59262 21940 59304 21996
rect 59164 21912 59304 21940
rect 59334 22236 59450 22264
rect 59334 22180 59364 22236
rect 59420 22180 59450 22236
rect 59334 22156 59450 22180
rect 59334 22100 59364 22156
rect 59420 22100 59450 22156
rect 59334 22076 59450 22100
rect 59334 22020 59364 22076
rect 59420 22020 59450 22076
rect 59334 21996 59450 22020
rect 59334 21940 59364 21996
rect 59420 21940 59450 21996
rect 59334 21912 59450 21940
rect 59642 22236 59758 22264
rect 59642 22180 59672 22236
rect 59728 22180 59758 22236
rect 59642 22156 59758 22180
rect 59642 22100 59672 22156
rect 59728 22100 59758 22156
rect 59642 22076 59758 22100
rect 59642 22020 59672 22076
rect 59728 22020 59758 22076
rect 59642 21996 59758 22020
rect 59642 21940 59672 21996
rect 59728 21940 59758 21996
rect 59642 21912 59758 21940
rect 59788 22236 59904 22264
rect 59788 22180 59818 22236
rect 59874 22180 59904 22236
rect 59788 22156 59904 22180
rect 59788 22100 59818 22156
rect 59874 22100 59904 22156
rect 59788 22076 59904 22100
rect 59788 22020 59818 22076
rect 59874 22020 59904 22076
rect 59788 21996 59904 22020
rect 59788 21940 59818 21996
rect 59874 21940 59904 21996
rect 59788 21912 59904 21940
rect 59934 22236 60110 22264
rect 59934 22180 59954 22236
rect 60010 22180 60034 22236
rect 60090 22180 60110 22236
rect 59934 22156 60110 22180
rect 59934 22100 59954 22156
rect 60010 22100 60034 22156
rect 60090 22100 60110 22156
rect 59934 22076 60110 22100
rect 59934 22020 59954 22076
rect 60010 22020 60034 22076
rect 60090 22020 60110 22076
rect 59934 21996 60110 22020
rect 59934 21940 59954 21996
rect 60010 21940 60034 21996
rect 60090 21940 60110 21996
rect 59934 21912 60110 21940
rect 62307 22236 62481 22264
rect 62307 22180 62326 22236
rect 62382 22180 62406 22236
rect 62462 22180 62481 22236
rect 62307 22156 62481 22180
rect 62307 22100 62326 22156
rect 62382 22100 62406 22156
rect 62462 22100 62481 22156
rect 62307 22076 62481 22100
rect 62307 22020 62326 22076
rect 62382 22020 62406 22076
rect 62462 22020 62481 22076
rect 62307 21996 62481 22020
rect 62307 21940 62326 21996
rect 62382 21940 62406 21996
rect 62462 21940 62481 21996
rect 62307 21912 62481 21940
rect 2020 14588 2124 14616
rect 2020 14532 2044 14588
rect 2100 14532 2124 14588
rect 2020 14508 2124 14532
rect 2020 14452 2044 14508
rect 2100 14452 2124 14508
rect 2020 14428 2124 14452
rect 2020 14372 2044 14428
rect 2100 14372 2124 14428
rect 2020 14348 2124 14372
rect 2020 14292 2044 14348
rect 2100 14292 2124 14348
rect 2020 14264 2124 14292
rect 5521 14588 5615 14616
rect 5521 14532 5540 14588
rect 5596 14532 5615 14588
rect 5521 14508 5615 14532
rect 5521 14452 5540 14508
rect 5596 14452 5615 14508
rect 5521 14428 5615 14452
rect 5521 14372 5540 14428
rect 5596 14372 5615 14428
rect 5521 14348 5615 14372
rect 5521 14292 5540 14348
rect 5596 14292 5615 14348
rect 5521 14264 5615 14292
rect 8411 14588 8505 14616
rect 8411 14532 8430 14588
rect 8486 14532 8505 14588
rect 8411 14508 8505 14532
rect 8411 14452 8430 14508
rect 8486 14452 8505 14508
rect 8411 14428 8505 14452
rect 8411 14372 8430 14428
rect 8486 14372 8505 14428
rect 8411 14348 8505 14372
rect 8411 14292 8430 14348
rect 8486 14292 8505 14348
rect 8411 14264 8505 14292
rect 11301 14588 11395 14616
rect 11301 14532 11320 14588
rect 11376 14532 11395 14588
rect 11301 14508 11395 14532
rect 11301 14452 11320 14508
rect 11376 14452 11395 14508
rect 11301 14428 11395 14452
rect 11301 14372 11320 14428
rect 11376 14372 11395 14428
rect 11301 14348 11395 14372
rect 11301 14292 11320 14348
rect 11376 14292 11395 14348
rect 11301 14264 11395 14292
rect 14191 14588 14285 14616
rect 14191 14532 14210 14588
rect 14266 14532 14285 14588
rect 14191 14508 14285 14532
rect 14191 14452 14210 14508
rect 14266 14452 14285 14508
rect 14191 14428 14285 14452
rect 14191 14372 14210 14428
rect 14266 14372 14285 14428
rect 14191 14348 14285 14372
rect 14191 14292 14210 14348
rect 14266 14292 14285 14348
rect 14191 14264 14285 14292
rect 17081 14588 17175 14616
rect 17081 14532 17100 14588
rect 17156 14532 17175 14588
rect 17081 14508 17175 14532
rect 17081 14452 17100 14508
rect 17156 14452 17175 14508
rect 17081 14428 17175 14452
rect 17081 14372 17100 14428
rect 17156 14372 17175 14428
rect 17081 14348 17175 14372
rect 17081 14292 17100 14348
rect 17156 14292 17175 14348
rect 17081 14264 17175 14292
rect 19971 14588 20065 14616
rect 19971 14532 19990 14588
rect 20046 14532 20065 14588
rect 19971 14508 20065 14532
rect 19971 14452 19990 14508
rect 20046 14452 20065 14508
rect 19971 14428 20065 14452
rect 19971 14372 19990 14428
rect 20046 14372 20065 14428
rect 19971 14348 20065 14372
rect 19971 14292 19990 14348
rect 20046 14292 20065 14348
rect 19971 14264 20065 14292
rect 22861 14588 22955 14616
rect 22861 14532 22880 14588
rect 22936 14532 22955 14588
rect 22861 14508 22955 14532
rect 22861 14452 22880 14508
rect 22936 14452 22955 14508
rect 22861 14428 22955 14452
rect 22861 14372 22880 14428
rect 22936 14372 22955 14428
rect 22861 14348 22955 14372
rect 22861 14292 22880 14348
rect 22936 14292 22955 14348
rect 22861 14264 22955 14292
rect 25751 14588 25845 14616
rect 25751 14532 25770 14588
rect 25826 14532 25845 14588
rect 25751 14508 25845 14532
rect 25751 14452 25770 14508
rect 25826 14452 25845 14508
rect 25751 14428 25845 14452
rect 25751 14372 25770 14428
rect 25826 14372 25845 14428
rect 25751 14348 25845 14372
rect 25751 14292 25770 14348
rect 25826 14292 25845 14348
rect 25751 14264 25845 14292
rect 28641 14588 28735 14616
rect 28641 14532 28660 14588
rect 28716 14532 28735 14588
rect 28641 14508 28735 14532
rect 28641 14452 28660 14508
rect 28716 14452 28735 14508
rect 28641 14428 28735 14452
rect 28641 14372 28660 14428
rect 28716 14372 28735 14428
rect 28641 14348 28735 14372
rect 28641 14292 28660 14348
rect 28716 14292 28735 14348
rect 28641 14264 28735 14292
rect 31531 14588 31625 14616
rect 31531 14532 31550 14588
rect 31606 14532 31625 14588
rect 31531 14508 31625 14532
rect 31531 14452 31550 14508
rect 31606 14452 31625 14508
rect 31531 14428 31625 14452
rect 31531 14372 31550 14428
rect 31606 14372 31625 14428
rect 31531 14348 31625 14372
rect 31531 14292 31550 14348
rect 31606 14292 31625 14348
rect 31531 14264 31625 14292
rect 34421 14588 34515 14616
rect 34421 14532 34440 14588
rect 34496 14532 34515 14588
rect 34421 14508 34515 14532
rect 34421 14452 34440 14508
rect 34496 14452 34515 14508
rect 34421 14428 34515 14452
rect 34421 14372 34440 14428
rect 34496 14372 34515 14428
rect 34421 14348 34515 14372
rect 34421 14292 34440 14348
rect 34496 14292 34515 14348
rect 34421 14264 34515 14292
rect 37311 14588 37405 14616
rect 37311 14532 37330 14588
rect 37386 14532 37405 14588
rect 37311 14508 37405 14532
rect 37311 14452 37330 14508
rect 37386 14452 37405 14508
rect 37311 14428 37405 14452
rect 37311 14372 37330 14428
rect 37386 14372 37405 14428
rect 37311 14348 37405 14372
rect 37311 14292 37330 14348
rect 37386 14292 37405 14348
rect 37311 14264 37405 14292
rect 40201 14588 40295 14616
rect 40201 14532 40220 14588
rect 40276 14532 40295 14588
rect 40201 14508 40295 14532
rect 40201 14452 40220 14508
rect 40276 14452 40295 14508
rect 40201 14428 40295 14452
rect 40201 14372 40220 14428
rect 40276 14372 40295 14428
rect 40201 14348 40295 14372
rect 40201 14292 40220 14348
rect 40276 14292 40295 14348
rect 40201 14264 40295 14292
rect 43091 14588 43185 14616
rect 43091 14532 43110 14588
rect 43166 14532 43185 14588
rect 43091 14508 43185 14532
rect 43091 14452 43110 14508
rect 43166 14452 43185 14508
rect 43091 14428 43185 14452
rect 43091 14372 43110 14428
rect 43166 14372 43185 14428
rect 43091 14348 43185 14372
rect 43091 14292 43110 14348
rect 43166 14292 43185 14348
rect 43091 14264 43185 14292
rect 45981 14588 46075 14616
rect 45981 14532 46000 14588
rect 46056 14532 46075 14588
rect 45981 14508 46075 14532
rect 45981 14452 46000 14508
rect 46056 14452 46075 14508
rect 45981 14428 46075 14452
rect 45981 14372 46000 14428
rect 46056 14372 46075 14428
rect 45981 14348 46075 14372
rect 45981 14292 46000 14348
rect 46056 14292 46075 14348
rect 45981 14264 46075 14292
rect 48989 14588 49083 14616
rect 48989 14532 49008 14588
rect 49064 14532 49083 14588
rect 48989 14508 49083 14532
rect 48989 14452 49008 14508
rect 49064 14452 49083 14508
rect 48989 14428 49083 14452
rect 48989 14372 49008 14428
rect 49064 14372 49083 14428
rect 48989 14348 49083 14372
rect 48989 14292 49008 14348
rect 49064 14292 49083 14348
rect 48989 14264 49083 14292
rect 52210 14588 52320 14616
rect 52210 14532 52237 14588
rect 52293 14532 52320 14588
rect 52210 14508 52320 14532
rect 52210 14452 52237 14508
rect 52293 14452 52320 14508
rect 52210 14428 52320 14452
rect 52210 14372 52237 14428
rect 52293 14372 52320 14428
rect 52210 14348 52320 14372
rect 52210 14292 52237 14348
rect 52293 14292 52320 14348
rect 52210 14264 52320 14292
rect 53602 14588 53730 14616
rect 53602 14532 53638 14588
rect 53694 14532 53730 14588
rect 53602 14508 53730 14532
rect 53602 14452 53638 14508
rect 53694 14452 53730 14508
rect 53602 14428 53730 14452
rect 53602 14372 53638 14428
rect 53694 14372 53730 14428
rect 53602 14348 53730 14372
rect 53602 14292 53638 14348
rect 53694 14292 53730 14348
rect 53602 14264 53730 14292
rect 53770 14588 53898 14616
rect 53770 14532 53806 14588
rect 53862 14532 53898 14588
rect 53770 14508 53898 14532
rect 53770 14452 53806 14508
rect 53862 14452 53898 14508
rect 53770 14428 53898 14452
rect 53770 14372 53806 14428
rect 53862 14372 53898 14428
rect 53770 14348 53898 14372
rect 53770 14292 53806 14348
rect 53862 14292 53898 14348
rect 53770 14264 53898 14292
rect 54514 14588 54642 14616
rect 54514 14532 54550 14588
rect 54606 14532 54642 14588
rect 54514 14508 54642 14532
rect 54514 14452 54550 14508
rect 54606 14452 54642 14508
rect 54514 14428 54642 14452
rect 54514 14372 54550 14428
rect 54606 14372 54642 14428
rect 54514 14348 54642 14372
rect 54514 14292 54550 14348
rect 54606 14292 54642 14348
rect 54514 14264 54642 14292
rect 54910 14588 55026 14616
rect 54910 14532 54940 14588
rect 54996 14532 55026 14588
rect 54910 14508 55026 14532
rect 54910 14452 54940 14508
rect 54996 14452 55026 14508
rect 54910 14428 55026 14452
rect 54910 14372 54940 14428
rect 54996 14372 55026 14428
rect 54910 14348 55026 14372
rect 54910 14292 54940 14348
rect 54996 14292 55026 14348
rect 54910 14264 55026 14292
rect 55620 14588 55748 14616
rect 55620 14532 55656 14588
rect 55712 14532 55748 14588
rect 55620 14508 55748 14532
rect 55620 14452 55656 14508
rect 55712 14452 55748 14508
rect 55620 14428 55748 14452
rect 55620 14372 55656 14428
rect 55712 14372 55748 14428
rect 55620 14348 55748 14372
rect 55620 14292 55656 14348
rect 55712 14292 55748 14348
rect 55620 14264 55748 14292
rect 56198 14588 56326 14616
rect 56198 14532 56234 14588
rect 56290 14532 56326 14588
rect 56198 14508 56326 14532
rect 56198 14452 56234 14508
rect 56290 14452 56326 14508
rect 56198 14428 56326 14452
rect 56198 14372 56234 14428
rect 56290 14372 56326 14428
rect 56198 14348 56326 14372
rect 56198 14292 56234 14348
rect 56290 14292 56326 14348
rect 56198 14264 56326 14292
rect 56649 14588 56765 14616
rect 56649 14532 56679 14588
rect 56735 14532 56765 14588
rect 56649 14508 56765 14532
rect 56649 14452 56679 14508
rect 56735 14452 56765 14508
rect 56649 14428 56765 14452
rect 56649 14372 56679 14428
rect 56735 14372 56765 14428
rect 56649 14348 56765 14372
rect 56649 14292 56679 14348
rect 56735 14292 56765 14348
rect 56649 14264 56765 14292
rect 56953 14588 57069 14616
rect 56953 14532 56983 14588
rect 57039 14532 57069 14588
rect 56953 14508 57069 14532
rect 56953 14452 56983 14508
rect 57039 14452 57069 14508
rect 56953 14428 57069 14452
rect 56953 14372 56983 14428
rect 57039 14372 57069 14428
rect 56953 14348 57069 14372
rect 56953 14292 56983 14348
rect 57039 14292 57069 14348
rect 56953 14264 57069 14292
rect 57795 14588 57911 14616
rect 57795 14532 57825 14588
rect 57881 14532 57911 14588
rect 57795 14508 57911 14532
rect 57795 14452 57825 14508
rect 57881 14452 57911 14508
rect 57795 14428 57911 14452
rect 57795 14372 57825 14428
rect 57881 14372 57911 14428
rect 57795 14348 57911 14372
rect 57795 14292 57825 14348
rect 57881 14292 57911 14348
rect 57795 14264 57911 14292
rect 58461 14588 58525 14616
rect 58461 14532 58465 14588
rect 58521 14532 58525 14588
rect 58461 14508 58525 14532
rect 58461 14452 58465 14508
rect 58521 14452 58525 14508
rect 58461 14428 58525 14452
rect 58461 14372 58465 14428
rect 58521 14372 58525 14428
rect 58461 14348 58525 14372
rect 58461 14292 58465 14348
rect 58521 14292 58525 14348
rect 58461 14264 58525 14292
rect 59018 14588 59134 14616
rect 59018 14532 59048 14588
rect 59104 14532 59134 14588
rect 59018 14508 59134 14532
rect 59018 14452 59048 14508
rect 59104 14452 59134 14508
rect 59018 14428 59134 14452
rect 59018 14372 59048 14428
rect 59104 14372 59134 14428
rect 59018 14348 59134 14372
rect 59018 14292 59048 14348
rect 59104 14292 59134 14348
rect 59018 14264 59134 14292
rect 60296 14588 60412 14616
rect 60296 14532 60326 14588
rect 60382 14532 60412 14588
rect 60296 14508 60412 14532
rect 60296 14452 60326 14508
rect 60382 14452 60412 14508
rect 60296 14428 60412 14452
rect 60296 14372 60326 14428
rect 60382 14372 60412 14428
rect 60296 14348 60412 14372
rect 60296 14292 60326 14348
rect 60382 14292 60412 14348
rect 60296 14264 60412 14292
rect 60454 14588 60570 14616
rect 60454 14532 60484 14588
rect 60540 14532 60570 14588
rect 60454 14508 60570 14532
rect 60454 14452 60484 14508
rect 60540 14452 60570 14508
rect 60454 14428 60570 14452
rect 60454 14372 60484 14428
rect 60540 14372 60570 14428
rect 60454 14348 60570 14372
rect 60454 14292 60484 14348
rect 60540 14292 60570 14348
rect 60454 14264 60570 14292
rect 62509 14588 62683 14616
rect 62509 14532 62528 14588
rect 62584 14532 62608 14588
rect 62664 14532 62683 14588
rect 62509 14508 62683 14532
rect 62509 14452 62528 14508
rect 62584 14452 62608 14508
rect 62664 14452 62683 14508
rect 62509 14428 62683 14452
rect 62509 14372 62528 14428
rect 62584 14372 62608 14428
rect 62664 14372 62683 14428
rect 62509 14348 62683 14372
rect 62509 14292 62528 14348
rect 62584 14292 62608 14348
rect 62664 14292 62683 14348
rect 62509 14264 62683 14292
rect 2152 12236 2352 12264
rect 2152 12180 2184 12236
rect 2240 12180 2264 12236
rect 2320 12180 2352 12236
rect 2152 12156 2352 12180
rect 2152 12100 2184 12156
rect 2240 12100 2264 12156
rect 2320 12100 2352 12156
rect 2152 12076 2352 12100
rect 2152 12020 2184 12076
rect 2240 12020 2264 12076
rect 2320 12020 2352 12076
rect 2152 11996 2352 12020
rect 2152 11940 2184 11996
rect 2240 11940 2264 11996
rect 2320 11940 2352 11996
rect 2152 11912 2352 11940
rect 5374 12236 5468 12264
rect 5374 12180 5393 12236
rect 5449 12180 5468 12236
rect 5374 12156 5468 12180
rect 5374 12100 5393 12156
rect 5449 12100 5468 12156
rect 5374 12076 5468 12100
rect 5374 12020 5393 12076
rect 5449 12020 5468 12076
rect 5374 11996 5468 12020
rect 5374 11940 5393 11996
rect 5449 11940 5468 11996
rect 5374 11912 5468 11940
rect 8264 12236 8358 12264
rect 8264 12180 8283 12236
rect 8339 12180 8358 12236
rect 8264 12156 8358 12180
rect 8264 12100 8283 12156
rect 8339 12100 8358 12156
rect 8264 12076 8358 12100
rect 8264 12020 8283 12076
rect 8339 12020 8358 12076
rect 8264 11996 8358 12020
rect 8264 11940 8283 11996
rect 8339 11940 8358 11996
rect 8264 11912 8358 11940
rect 11154 12236 11248 12264
rect 11154 12180 11173 12236
rect 11229 12180 11248 12236
rect 11154 12156 11248 12180
rect 11154 12100 11173 12156
rect 11229 12100 11248 12156
rect 11154 12076 11248 12100
rect 11154 12020 11173 12076
rect 11229 12020 11248 12076
rect 11154 11996 11248 12020
rect 11154 11940 11173 11996
rect 11229 11940 11248 11996
rect 11154 11912 11248 11940
rect 14044 12236 14138 12264
rect 14044 12180 14063 12236
rect 14119 12180 14138 12236
rect 14044 12156 14138 12180
rect 14044 12100 14063 12156
rect 14119 12100 14138 12156
rect 14044 12076 14138 12100
rect 14044 12020 14063 12076
rect 14119 12020 14138 12076
rect 14044 11996 14138 12020
rect 14044 11940 14063 11996
rect 14119 11940 14138 11996
rect 14044 11912 14138 11940
rect 16934 12236 17028 12264
rect 16934 12180 16953 12236
rect 17009 12180 17028 12236
rect 16934 12156 17028 12180
rect 16934 12100 16953 12156
rect 17009 12100 17028 12156
rect 16934 12076 17028 12100
rect 16934 12020 16953 12076
rect 17009 12020 17028 12076
rect 16934 11996 17028 12020
rect 16934 11940 16953 11996
rect 17009 11940 17028 11996
rect 16934 11912 17028 11940
rect 19824 12236 19918 12264
rect 19824 12180 19843 12236
rect 19899 12180 19918 12236
rect 19824 12156 19918 12180
rect 19824 12100 19843 12156
rect 19899 12100 19918 12156
rect 19824 12076 19918 12100
rect 19824 12020 19843 12076
rect 19899 12020 19918 12076
rect 19824 11996 19918 12020
rect 19824 11940 19843 11996
rect 19899 11940 19918 11996
rect 19824 11912 19918 11940
rect 22714 12236 22808 12264
rect 22714 12180 22733 12236
rect 22789 12180 22808 12236
rect 22714 12156 22808 12180
rect 22714 12100 22733 12156
rect 22789 12100 22808 12156
rect 22714 12076 22808 12100
rect 22714 12020 22733 12076
rect 22789 12020 22808 12076
rect 22714 11996 22808 12020
rect 22714 11940 22733 11996
rect 22789 11940 22808 11996
rect 22714 11912 22808 11940
rect 25604 12236 25698 12264
rect 25604 12180 25623 12236
rect 25679 12180 25698 12236
rect 25604 12156 25698 12180
rect 25604 12100 25623 12156
rect 25679 12100 25698 12156
rect 25604 12076 25698 12100
rect 25604 12020 25623 12076
rect 25679 12020 25698 12076
rect 25604 11996 25698 12020
rect 25604 11940 25623 11996
rect 25679 11940 25698 11996
rect 25604 11912 25698 11940
rect 28494 12236 28588 12264
rect 28494 12180 28513 12236
rect 28569 12180 28588 12236
rect 28494 12156 28588 12180
rect 28494 12100 28513 12156
rect 28569 12100 28588 12156
rect 28494 12076 28588 12100
rect 28494 12020 28513 12076
rect 28569 12020 28588 12076
rect 28494 11996 28588 12020
rect 28494 11940 28513 11996
rect 28569 11940 28588 11996
rect 28494 11912 28588 11940
rect 31384 12236 31478 12264
rect 31384 12180 31403 12236
rect 31459 12180 31478 12236
rect 31384 12156 31478 12180
rect 31384 12100 31403 12156
rect 31459 12100 31478 12156
rect 31384 12076 31478 12100
rect 31384 12020 31403 12076
rect 31459 12020 31478 12076
rect 31384 11996 31478 12020
rect 31384 11940 31403 11996
rect 31459 11940 31478 11996
rect 31384 11912 31478 11940
rect 34274 12236 34368 12264
rect 34274 12180 34293 12236
rect 34349 12180 34368 12236
rect 34274 12156 34368 12180
rect 34274 12100 34293 12156
rect 34349 12100 34368 12156
rect 34274 12076 34368 12100
rect 34274 12020 34293 12076
rect 34349 12020 34368 12076
rect 34274 11996 34368 12020
rect 34274 11940 34293 11996
rect 34349 11940 34368 11996
rect 34274 11912 34368 11940
rect 37164 12236 37258 12264
rect 37164 12180 37183 12236
rect 37239 12180 37258 12236
rect 37164 12156 37258 12180
rect 37164 12100 37183 12156
rect 37239 12100 37258 12156
rect 37164 12076 37258 12100
rect 37164 12020 37183 12076
rect 37239 12020 37258 12076
rect 37164 11996 37258 12020
rect 37164 11940 37183 11996
rect 37239 11940 37258 11996
rect 37164 11912 37258 11940
rect 40054 12236 40148 12264
rect 40054 12180 40073 12236
rect 40129 12180 40148 12236
rect 40054 12156 40148 12180
rect 40054 12100 40073 12156
rect 40129 12100 40148 12156
rect 40054 12076 40148 12100
rect 40054 12020 40073 12076
rect 40129 12020 40148 12076
rect 40054 11996 40148 12020
rect 40054 11940 40073 11996
rect 40129 11940 40148 11996
rect 40054 11912 40148 11940
rect 42944 12236 43038 12264
rect 42944 12180 42963 12236
rect 43019 12180 43038 12236
rect 42944 12156 43038 12180
rect 42944 12100 42963 12156
rect 43019 12100 43038 12156
rect 42944 12076 43038 12100
rect 42944 12020 42963 12076
rect 43019 12020 43038 12076
rect 42944 11996 43038 12020
rect 42944 11940 42963 11996
rect 43019 11940 43038 11996
rect 42944 11912 43038 11940
rect 45834 12236 45928 12264
rect 45834 12180 45853 12236
rect 45909 12180 45928 12236
rect 45834 12156 45928 12180
rect 45834 12100 45853 12156
rect 45909 12100 45928 12156
rect 45834 12076 45928 12100
rect 45834 12020 45853 12076
rect 45909 12020 45928 12076
rect 45834 11996 45928 12020
rect 45834 11940 45853 11996
rect 45909 11940 45928 11996
rect 45834 11912 45928 11940
rect 48781 12236 48875 12264
rect 48781 12180 48800 12236
rect 48856 12180 48875 12236
rect 48781 12156 48875 12180
rect 48781 12100 48800 12156
rect 48856 12100 48875 12156
rect 48781 12076 48875 12100
rect 48781 12020 48800 12076
rect 48856 12020 48875 12076
rect 48781 11996 48875 12020
rect 48781 11940 48800 11996
rect 48856 11940 48875 11996
rect 48781 11912 48875 11940
rect 49630 12236 49830 12264
rect 49630 12180 49662 12236
rect 49718 12180 49742 12236
rect 49798 12180 49830 12236
rect 49630 12156 49830 12180
rect 49630 12100 49662 12156
rect 49718 12100 49742 12156
rect 49798 12100 49830 12156
rect 49630 12076 49830 12100
rect 49630 12020 49662 12076
rect 49718 12020 49742 12076
rect 49798 12020 49830 12076
rect 49630 11996 49830 12020
rect 49630 11940 49662 11996
rect 49718 11940 49742 11996
rect 49798 11940 49830 11996
rect 49630 11912 49830 11940
rect 52920 12236 53048 12264
rect 52920 12180 52956 12236
rect 53012 12180 53048 12236
rect 52920 12156 53048 12180
rect 52920 12100 52956 12156
rect 53012 12100 53048 12156
rect 52920 12076 53048 12100
rect 52920 12020 52956 12076
rect 53012 12020 53048 12076
rect 52920 11996 53048 12020
rect 52920 11940 52956 11996
rect 53012 11940 53048 11996
rect 52920 11912 53048 11940
rect 53078 12236 53206 12264
rect 53078 12180 53114 12236
rect 53170 12180 53206 12236
rect 53078 12156 53206 12180
rect 53078 12100 53114 12156
rect 53170 12100 53206 12156
rect 53078 12076 53206 12100
rect 53078 12020 53114 12076
rect 53170 12020 53206 12076
rect 53078 11996 53206 12020
rect 53078 11940 53114 11996
rect 53170 11940 53206 11996
rect 53078 11912 53206 11940
rect 53434 12236 53562 12264
rect 53434 12180 53470 12236
rect 53526 12180 53562 12236
rect 53434 12156 53562 12180
rect 53434 12100 53470 12156
rect 53526 12100 53562 12156
rect 53434 12076 53562 12100
rect 53434 12020 53470 12076
rect 53526 12020 53562 12076
rect 53434 11996 53562 12020
rect 53434 11940 53470 11996
rect 53526 11940 53562 11996
rect 53434 11912 53562 11940
rect 54752 12236 54880 12264
rect 54752 12180 54788 12236
rect 54844 12180 54880 12236
rect 54752 12156 54880 12180
rect 54752 12100 54788 12156
rect 54844 12100 54880 12156
rect 54752 12076 54880 12100
rect 54752 12020 54788 12076
rect 54844 12020 54880 12076
rect 54752 11996 54880 12020
rect 54752 11940 54788 11996
rect 54844 11940 54880 11996
rect 54752 11912 54880 11940
rect 55345 12236 55473 12264
rect 55345 12180 55381 12236
rect 55437 12180 55473 12236
rect 55345 12156 55473 12180
rect 55345 12100 55381 12156
rect 55437 12100 55473 12156
rect 55345 12076 55473 12100
rect 55345 12020 55381 12076
rect 55437 12020 55473 12076
rect 55345 11996 55473 12020
rect 55345 11940 55381 11996
rect 55437 11940 55473 11996
rect 55345 11912 55473 11940
rect 56491 12236 56619 12264
rect 56491 12180 56527 12236
rect 56583 12180 56619 12236
rect 56491 12156 56619 12180
rect 56491 12100 56527 12156
rect 56583 12100 56619 12156
rect 56491 12076 56619 12100
rect 56491 12020 56527 12076
rect 56583 12020 56619 12076
rect 56491 11996 56619 12020
rect 56491 11940 56527 11996
rect 56583 11940 56619 11996
rect 56491 11912 56619 11940
rect 57941 12236 58121 12264
rect 57941 12180 57963 12236
rect 58019 12180 58043 12236
rect 58099 12180 58121 12236
rect 57941 12156 58121 12180
rect 57941 12100 57963 12156
rect 58019 12100 58043 12156
rect 58099 12100 58121 12156
rect 57941 12076 58121 12100
rect 57941 12020 57963 12076
rect 58019 12020 58043 12076
rect 58099 12020 58121 12076
rect 57941 11996 58121 12020
rect 57941 11940 57963 11996
rect 58019 11940 58043 11996
rect 58099 11940 58121 11996
rect 57941 11912 58121 11940
rect 59164 12236 59304 12264
rect 59164 12180 59206 12236
rect 59262 12180 59304 12236
rect 59164 12156 59304 12180
rect 59164 12100 59206 12156
rect 59262 12100 59304 12156
rect 59164 12076 59304 12100
rect 59164 12020 59206 12076
rect 59262 12020 59304 12076
rect 59164 11996 59304 12020
rect 59164 11940 59206 11996
rect 59262 11940 59304 11996
rect 59164 11912 59304 11940
rect 59334 12236 59450 12264
rect 59334 12180 59364 12236
rect 59420 12180 59450 12236
rect 59334 12156 59450 12180
rect 59334 12100 59364 12156
rect 59420 12100 59450 12156
rect 59334 12076 59450 12100
rect 59334 12020 59364 12076
rect 59420 12020 59450 12076
rect 59334 11996 59450 12020
rect 59334 11940 59364 11996
rect 59420 11940 59450 11996
rect 59334 11912 59450 11940
rect 59642 12236 59758 12264
rect 59642 12180 59672 12236
rect 59728 12180 59758 12236
rect 59642 12156 59758 12180
rect 59642 12100 59672 12156
rect 59728 12100 59758 12156
rect 59642 12076 59758 12100
rect 59642 12020 59672 12076
rect 59728 12020 59758 12076
rect 59642 11996 59758 12020
rect 59642 11940 59672 11996
rect 59728 11940 59758 11996
rect 59642 11912 59758 11940
rect 59788 12236 59904 12264
rect 59788 12180 59818 12236
rect 59874 12180 59904 12236
rect 59788 12156 59904 12180
rect 59788 12100 59818 12156
rect 59874 12100 59904 12156
rect 59788 12076 59904 12100
rect 59788 12020 59818 12076
rect 59874 12020 59904 12076
rect 59788 11996 59904 12020
rect 59788 11940 59818 11996
rect 59874 11940 59904 11996
rect 59788 11912 59904 11940
rect 59934 12236 60110 12264
rect 59934 12180 59954 12236
rect 60010 12180 60034 12236
rect 60090 12180 60110 12236
rect 59934 12156 60110 12180
rect 59934 12100 59954 12156
rect 60010 12100 60034 12156
rect 60090 12100 60110 12156
rect 59934 12076 60110 12100
rect 59934 12020 59954 12076
rect 60010 12020 60034 12076
rect 60090 12020 60110 12076
rect 59934 11996 60110 12020
rect 59934 11940 59954 11996
rect 60010 11940 60034 11996
rect 60090 11940 60110 11996
rect 59934 11912 60110 11940
rect 62307 12236 62481 12264
rect 62307 12180 62326 12236
rect 62382 12180 62406 12236
rect 62462 12180 62481 12236
rect 62307 12156 62481 12180
rect 62307 12100 62326 12156
rect 62382 12100 62406 12156
rect 62462 12100 62481 12156
rect 62307 12076 62481 12100
rect 62307 12020 62326 12076
rect 62382 12020 62406 12076
rect 62462 12020 62481 12076
rect 62307 11996 62481 12020
rect 62307 11940 62326 11996
rect 62382 11940 62406 11996
rect 62462 11940 62481 11996
rect 62307 11912 62481 11940
rect 63420 11234 63448 38878
rect 63512 11422 63540 61172
rect 63500 11416 63552 11422
rect 63500 11358 63552 11364
rect 63604 11354 63632 63038
rect 63684 56636 63736 56642
rect 63684 56578 63736 56584
rect 63592 11348 63644 11354
rect 63592 11290 63644 11296
rect 63420 11206 63632 11234
rect 63408 11144 63460 11150
rect 63408 11086 63460 11092
rect 59196 7886 59224 8024
rect 59184 7880 59236 7886
rect 59184 7822 59236 7828
rect 59572 7818 59600 8024
rect 63224 7880 63276 7886
rect 63224 7822 63276 7828
rect 47308 7812 47360 7818
rect 47308 7754 47360 7760
rect 55772 7812 55824 7818
rect 55772 7754 55824 7760
rect 59560 7812 59612 7818
rect 59560 7754 59612 7760
rect 44824 7744 44876 7750
rect 44824 7686 44876 7692
rect 33048 7608 33100 7614
rect 33048 7550 33100 7556
rect 1836 4922 2188 5944
rect 1836 4870 1858 4922
rect 1910 4870 1922 4922
rect 1974 4870 1986 4922
rect 2038 4870 2050 4922
rect 2102 4870 2114 4922
rect 2166 4870 2188 4922
rect 1836 3834 2188 4870
rect 1836 3782 1858 3834
rect 1910 3782 1922 3834
rect 1974 3782 1986 3834
rect 2038 3782 2050 3834
rect 2102 3782 2114 3834
rect 2166 3782 2188 3834
rect 1836 2746 2188 3782
rect 1836 2694 1858 2746
rect 1910 2694 1922 2746
rect 1974 2694 1986 2746
rect 2038 2694 2050 2746
rect 2102 2694 2114 2746
rect 2166 2694 2188 2746
rect 1836 2236 2188 2694
rect 1836 2180 1864 2236
rect 1920 2180 1944 2236
rect 2000 2180 2024 2236
rect 2080 2180 2104 2236
rect 2160 2180 2188 2236
rect 1836 2156 2188 2180
rect 1836 2100 1864 2156
rect 1920 2100 1944 2156
rect 2000 2100 2024 2156
rect 2080 2100 2104 2156
rect 2160 2100 2188 2156
rect 1836 2076 2188 2100
rect 1836 2020 1864 2076
rect 1920 2020 1944 2076
rect 2000 2020 2024 2076
rect 2080 2020 2104 2076
rect 2160 2020 2188 2076
rect 1836 1996 2188 2020
rect 1836 1940 1864 1996
rect 1920 1940 1944 1996
rect 2000 1940 2024 1996
rect 2080 1940 2104 1996
rect 2160 1940 2188 1996
rect 1836 1658 2188 1940
rect 1836 1606 1858 1658
rect 1910 1606 1922 1658
rect 1974 1606 1986 1658
rect 2038 1606 2050 1658
rect 2102 1606 2114 1658
rect 2166 1606 2188 1658
rect 1836 1040 2188 1606
rect 4188 5466 4540 5972
rect 4188 5414 4210 5466
rect 4262 5414 4274 5466
rect 4326 5414 4338 5466
rect 4390 5414 4402 5466
rect 4454 5414 4466 5466
rect 4518 5414 4540 5466
rect 4188 4588 4540 5414
rect 4188 4532 4216 4588
rect 4272 4532 4296 4588
rect 4352 4532 4376 4588
rect 4432 4532 4456 4588
rect 4512 4532 4540 4588
rect 4188 4508 4540 4532
rect 4188 4452 4216 4508
rect 4272 4452 4296 4508
rect 4352 4452 4376 4508
rect 4432 4452 4456 4508
rect 4512 4452 4540 4508
rect 4188 4428 4540 4452
rect 4188 4378 4216 4428
rect 4272 4378 4296 4428
rect 4352 4378 4376 4428
rect 4432 4378 4456 4428
rect 4512 4378 4540 4428
rect 4188 4326 4210 4378
rect 4272 4372 4274 4378
rect 4454 4372 4456 4378
rect 4262 4348 4274 4372
rect 4326 4348 4338 4372
rect 4390 4348 4402 4372
rect 4454 4348 4466 4372
rect 4272 4326 4274 4348
rect 4454 4326 4456 4348
rect 4518 4326 4540 4378
rect 4188 4292 4216 4326
rect 4272 4292 4296 4326
rect 4352 4292 4376 4326
rect 4432 4292 4456 4326
rect 4512 4292 4540 4326
rect 4188 3290 4540 4292
rect 4188 3238 4210 3290
rect 4262 3238 4274 3290
rect 4326 3238 4338 3290
rect 4390 3238 4402 3290
rect 4454 3238 4466 3290
rect 4518 3238 4540 3290
rect 4188 2202 4540 3238
rect 4188 2150 4210 2202
rect 4262 2150 4274 2202
rect 4326 2150 4338 2202
rect 4390 2150 4402 2202
rect 4454 2150 4466 2202
rect 4518 2150 4540 2202
rect 4188 1114 4540 2150
rect 4188 1062 4210 1114
rect 4262 1062 4274 1114
rect 4326 1062 4338 1114
rect 4390 1062 4402 1114
rect 4454 1062 4466 1114
rect 4518 1062 4540 1114
rect 4188 1040 4540 1062
rect 11836 4922 12188 5972
rect 11836 4870 11858 4922
rect 11910 4870 11922 4922
rect 11974 4870 11986 4922
rect 12038 4870 12050 4922
rect 12102 4870 12114 4922
rect 12166 4870 12188 4922
rect 11836 3834 12188 4870
rect 11836 3782 11858 3834
rect 11910 3782 11922 3834
rect 11974 3782 11986 3834
rect 12038 3782 12050 3834
rect 12102 3782 12114 3834
rect 12166 3782 12188 3834
rect 11836 2746 12188 3782
rect 11836 2694 11858 2746
rect 11910 2694 11922 2746
rect 11974 2694 11986 2746
rect 12038 2694 12050 2746
rect 12102 2694 12114 2746
rect 12166 2694 12188 2746
rect 11836 2236 12188 2694
rect 11836 2180 11864 2236
rect 11920 2180 11944 2236
rect 12000 2180 12024 2236
rect 12080 2180 12104 2236
rect 12160 2180 12188 2236
rect 11836 2156 12188 2180
rect 11836 2100 11864 2156
rect 11920 2100 11944 2156
rect 12000 2100 12024 2156
rect 12080 2100 12104 2156
rect 12160 2100 12188 2156
rect 11836 2076 12188 2100
rect 11836 2020 11864 2076
rect 11920 2020 11944 2076
rect 12000 2020 12024 2076
rect 12080 2020 12104 2076
rect 12160 2020 12188 2076
rect 11836 1996 12188 2020
rect 11836 1940 11864 1996
rect 11920 1940 11944 1996
rect 12000 1940 12024 1996
rect 12080 1940 12104 1996
rect 12160 1940 12188 1996
rect 11836 1658 12188 1940
rect 11836 1606 11858 1658
rect 11910 1606 11922 1658
rect 11974 1606 11986 1658
rect 12038 1606 12050 1658
rect 12102 1606 12114 1658
rect 12166 1606 12188 1658
rect 11836 1040 12188 1606
rect 14188 5466 14540 5972
rect 14188 5414 14210 5466
rect 14262 5414 14274 5466
rect 14326 5414 14338 5466
rect 14390 5414 14402 5466
rect 14454 5414 14466 5466
rect 14518 5414 14540 5466
rect 14188 4588 14540 5414
rect 14188 4532 14216 4588
rect 14272 4532 14296 4588
rect 14352 4532 14376 4588
rect 14432 4532 14456 4588
rect 14512 4532 14540 4588
rect 14188 4508 14540 4532
rect 14188 4452 14216 4508
rect 14272 4452 14296 4508
rect 14352 4452 14376 4508
rect 14432 4452 14456 4508
rect 14512 4452 14540 4508
rect 14188 4428 14540 4452
rect 14188 4378 14216 4428
rect 14272 4378 14296 4428
rect 14352 4378 14376 4428
rect 14432 4378 14456 4428
rect 14512 4378 14540 4428
rect 14188 4326 14210 4378
rect 14272 4372 14274 4378
rect 14454 4372 14456 4378
rect 14262 4348 14274 4372
rect 14326 4348 14338 4372
rect 14390 4348 14402 4372
rect 14454 4348 14466 4372
rect 14272 4326 14274 4348
rect 14454 4326 14456 4348
rect 14518 4326 14540 4378
rect 14188 4292 14216 4326
rect 14272 4292 14296 4326
rect 14352 4292 14376 4326
rect 14432 4292 14456 4326
rect 14512 4292 14540 4326
rect 14188 3290 14540 4292
rect 14188 3238 14210 3290
rect 14262 3238 14274 3290
rect 14326 3238 14338 3290
rect 14390 3238 14402 3290
rect 14454 3238 14466 3290
rect 14518 3238 14540 3290
rect 14188 2202 14540 3238
rect 21836 4922 22188 5972
rect 24188 5466 24540 5972
rect 28908 5704 28960 5710
rect 28908 5646 28960 5652
rect 29552 5704 29604 5710
rect 29552 5646 29604 5652
rect 30380 5704 30432 5710
rect 30380 5646 30432 5652
rect 30748 5704 30800 5710
rect 30748 5646 30800 5652
rect 31392 5704 31444 5710
rect 31392 5646 31444 5652
rect 24188 5414 24210 5466
rect 24262 5414 24274 5466
rect 24326 5414 24338 5466
rect 24390 5414 24402 5466
rect 24454 5414 24466 5466
rect 24518 5414 24540 5466
rect 23572 5092 23624 5098
rect 23572 5034 23624 5040
rect 21836 4870 21858 4922
rect 21910 4870 21922 4922
rect 21974 4870 21986 4922
rect 22038 4870 22050 4922
rect 22102 4870 22114 4922
rect 22166 4870 22188 4922
rect 21836 3834 22188 4870
rect 23480 4480 23532 4486
rect 23480 4422 23532 4428
rect 21836 3782 21858 3834
rect 21910 3782 21922 3834
rect 21974 3782 21986 3834
rect 22038 3782 22050 3834
rect 22102 3782 22114 3834
rect 22166 3782 22188 3834
rect 20996 2916 21048 2922
rect 20996 2858 21048 2864
rect 14188 2150 14210 2202
rect 14262 2150 14274 2202
rect 14326 2150 14338 2202
rect 14390 2150 14402 2202
rect 14454 2150 14466 2202
rect 14518 2150 14540 2202
rect 14188 1114 14540 2150
rect 21008 1358 21036 2858
rect 21836 2746 22188 3782
rect 23018 3360 23074 3369
rect 23018 3295 23074 3304
rect 22376 2984 22428 2990
rect 22376 2926 22428 2932
rect 22284 2848 22336 2854
rect 22284 2790 22336 2796
rect 21836 2694 21858 2746
rect 21910 2694 21922 2746
rect 21974 2694 21986 2746
rect 22038 2694 22050 2746
rect 22102 2694 22114 2746
rect 22166 2694 22188 2746
rect 21836 2236 22188 2694
rect 21836 2180 21864 2236
rect 21920 2180 21944 2236
rect 22000 2180 22024 2236
rect 22080 2180 22104 2236
rect 22160 2180 22188 2236
rect 21836 2156 22188 2180
rect 21836 2100 21864 2156
rect 21920 2100 21944 2156
rect 22000 2100 22024 2156
rect 22080 2100 22104 2156
rect 22160 2100 22188 2156
rect 21836 2076 22188 2100
rect 21836 2020 21864 2076
rect 21920 2020 21944 2076
rect 22000 2020 22024 2076
rect 22080 2020 22104 2076
rect 22160 2020 22188 2076
rect 21836 1996 22188 2020
rect 21836 1940 21864 1996
rect 21920 1940 21944 1996
rect 22000 1940 22024 1996
rect 22080 1940 22104 1996
rect 22160 1940 22188 1996
rect 21836 1658 22188 1940
rect 21836 1606 21858 1658
rect 21910 1606 21922 1658
rect 21974 1606 21986 1658
rect 22038 1606 22050 1658
rect 22102 1606 22114 1658
rect 22166 1606 22188 1658
rect 20996 1352 21048 1358
rect 20996 1294 21048 1300
rect 21732 1352 21784 1358
rect 21732 1294 21784 1300
rect 20812 1216 20864 1222
rect 20812 1158 20864 1164
rect 21548 1216 21600 1222
rect 21548 1158 21600 1164
rect 14188 1062 14210 1114
rect 14262 1062 14274 1114
rect 14326 1062 14338 1114
rect 14390 1062 14402 1114
rect 14454 1062 14466 1114
rect 14518 1062 14540 1114
rect 14188 1040 14540 1062
rect 20824 950 20852 1158
rect 20812 944 20864 950
rect 20812 886 20864 892
rect 21560 814 21588 1158
rect 21744 1018 21772 1294
rect 21836 1040 22188 1606
rect 22296 1222 22324 2790
rect 22388 2106 22416 2926
rect 22376 2100 22428 2106
rect 22376 2042 22428 2048
rect 22836 1760 22888 1766
rect 22836 1702 22888 1708
rect 22848 1426 22876 1702
rect 22376 1420 22428 1426
rect 22376 1362 22428 1368
rect 22836 1420 22888 1426
rect 22836 1362 22888 1368
rect 22284 1216 22336 1222
rect 22284 1158 22336 1164
rect 21732 1012 21784 1018
rect 21732 954 21784 960
rect 22388 882 22416 1362
rect 22652 1216 22704 1222
rect 22652 1158 22704 1164
rect 22376 876 22428 882
rect 22376 818 22428 824
rect 21548 808 21600 814
rect 21548 750 21600 756
rect 22664 746 22692 1158
rect 23032 800 23060 3295
rect 23112 2984 23164 2990
rect 23112 2926 23164 2932
rect 23124 2650 23152 2926
rect 23492 2854 23520 4422
rect 23584 2922 23612 5034
rect 24188 4588 24540 5414
rect 25044 5160 25096 5166
rect 25044 5102 25096 5108
rect 26148 5160 26200 5166
rect 26148 5102 26200 5108
rect 28356 5160 28408 5166
rect 28356 5102 28408 5108
rect 24188 4532 24216 4588
rect 24272 4532 24296 4588
rect 24352 4532 24376 4588
rect 24432 4532 24456 4588
rect 24512 4532 24540 4588
rect 24860 4616 24912 4622
rect 24860 4558 24912 4564
rect 24188 4508 24540 4532
rect 24188 4452 24216 4508
rect 24272 4452 24296 4508
rect 24352 4452 24376 4508
rect 24432 4452 24456 4508
rect 24512 4452 24540 4508
rect 24188 4428 24540 4452
rect 24188 4378 24216 4428
rect 24272 4378 24296 4428
rect 24352 4378 24376 4428
rect 24432 4378 24456 4428
rect 24512 4378 24540 4428
rect 24188 4326 24210 4378
rect 24272 4372 24274 4378
rect 24454 4372 24456 4378
rect 24262 4348 24274 4372
rect 24326 4348 24338 4372
rect 24390 4348 24402 4372
rect 24454 4348 24466 4372
rect 24272 4326 24274 4348
rect 24454 4326 24456 4348
rect 24518 4326 24540 4378
rect 24188 4292 24216 4326
rect 24272 4292 24296 4326
rect 24352 4292 24376 4326
rect 24432 4292 24456 4326
rect 24512 4292 24540 4326
rect 23664 3528 23716 3534
rect 23664 3470 23716 3476
rect 23572 2916 23624 2922
rect 23572 2858 23624 2864
rect 23480 2848 23532 2854
rect 23480 2790 23532 2796
rect 23112 2644 23164 2650
rect 23112 2586 23164 2592
rect 23480 2304 23532 2310
rect 23480 2246 23532 2252
rect 23492 1970 23520 2246
rect 23480 1964 23532 1970
rect 23480 1906 23532 1912
rect 23572 1896 23624 1902
rect 23572 1838 23624 1844
rect 23584 1562 23612 1838
rect 23572 1556 23624 1562
rect 23572 1498 23624 1504
rect 23388 1216 23440 1222
rect 23388 1158 23440 1164
rect 23400 1018 23428 1158
rect 23296 1012 23348 1018
rect 23296 954 23348 960
rect 23388 1012 23440 1018
rect 23388 954 23440 960
rect 23308 898 23336 954
rect 23676 950 23704 3470
rect 24032 3392 24084 3398
rect 24032 3334 24084 3340
rect 23848 2984 23900 2990
rect 23848 2926 23900 2932
rect 23860 2650 23888 2926
rect 23848 2644 23900 2650
rect 23848 2586 23900 2592
rect 24044 2582 24072 3334
rect 24188 3290 24540 4292
rect 24584 4072 24636 4078
rect 24584 4014 24636 4020
rect 24188 3238 24210 3290
rect 24262 3238 24274 3290
rect 24326 3238 24338 3290
rect 24390 3238 24402 3290
rect 24454 3238 24466 3290
rect 24518 3238 24540 3290
rect 24032 2576 24084 2582
rect 24032 2518 24084 2524
rect 24032 2440 24084 2446
rect 24032 2382 24084 2388
rect 24044 1902 24072 2382
rect 24188 2202 24540 3238
rect 24596 3194 24624 4014
rect 24584 3188 24636 3194
rect 24584 3130 24636 3136
rect 24584 2848 24636 2854
rect 24872 2802 24900 4558
rect 24952 3392 25004 3398
rect 24952 3334 25004 3340
rect 24584 2790 24636 2796
rect 24596 2378 24624 2790
rect 24780 2774 24900 2802
rect 24584 2372 24636 2378
rect 24584 2314 24636 2320
rect 24188 2150 24210 2202
rect 24262 2150 24274 2202
rect 24326 2150 24338 2202
rect 24390 2150 24402 2202
rect 24454 2150 24466 2202
rect 24518 2150 24540 2202
rect 24032 1896 24084 1902
rect 24032 1838 24084 1844
rect 23940 1284 23992 1290
rect 23940 1226 23992 1232
rect 23664 944 23716 950
rect 23308 870 23520 898
rect 23664 886 23716 892
rect 23492 800 23520 870
rect 23952 800 23980 1226
rect 24188 1114 24540 2150
rect 24188 1062 24210 1114
rect 24262 1062 24274 1114
rect 24326 1062 24338 1114
rect 24390 1062 24402 1114
rect 24454 1062 24466 1114
rect 24518 1062 24540 1114
rect 24188 1040 24540 1062
rect 24412 870 24532 898
rect 24412 800 24440 870
rect 22652 740 22704 746
rect 22652 682 22704 688
rect 23018 0 23074 800
rect 23478 0 23534 800
rect 23938 0 23994 800
rect 24398 0 24454 800
rect 24504 762 24532 870
rect 24780 762 24808 2774
rect 24964 2106 24992 3334
rect 25056 3058 25084 5102
rect 26160 4826 26188 5102
rect 26700 5024 26752 5030
rect 26700 4966 26752 4972
rect 27896 5024 27948 5030
rect 27896 4966 27948 4972
rect 26148 4820 26200 4826
rect 26148 4762 26200 4768
rect 26332 4684 26384 4690
rect 26332 4626 26384 4632
rect 26240 4616 26292 4622
rect 26240 4558 26292 4564
rect 25136 4072 25188 4078
rect 25136 4014 25188 4020
rect 25964 4072 26016 4078
rect 25964 4014 26016 4020
rect 25044 3052 25096 3058
rect 25044 2994 25096 3000
rect 24952 2100 25004 2106
rect 24952 2042 25004 2048
rect 24860 1760 24912 1766
rect 25148 1714 25176 4014
rect 25228 3936 25280 3942
rect 25228 3878 25280 3884
rect 25320 3936 25372 3942
rect 25320 3878 25372 3884
rect 25240 1970 25268 3878
rect 25332 3534 25360 3878
rect 25320 3528 25372 3534
rect 25320 3470 25372 3476
rect 25976 3126 26004 4014
rect 26056 3936 26108 3942
rect 26056 3878 26108 3884
rect 25964 3120 26016 3126
rect 25964 3062 26016 3068
rect 25320 2984 25372 2990
rect 25320 2926 25372 2932
rect 25332 2310 25360 2926
rect 25412 2848 25464 2854
rect 25412 2790 25464 2796
rect 25424 2446 25452 2790
rect 25412 2440 25464 2446
rect 25412 2382 25464 2388
rect 25320 2304 25372 2310
rect 25320 2246 25372 2252
rect 25228 1964 25280 1970
rect 25228 1906 25280 1912
rect 25320 1896 25372 1902
rect 25320 1838 25372 1844
rect 25596 1896 25648 1902
rect 25596 1838 25648 1844
rect 24860 1702 24912 1708
rect 24872 800 24900 1702
rect 25056 1686 25176 1714
rect 25056 814 25084 1686
rect 25136 1352 25188 1358
rect 25136 1294 25188 1300
rect 25148 814 25176 1294
rect 25044 808 25096 814
rect 24504 734 24808 762
rect 24858 0 24914 800
rect 25044 750 25096 756
rect 25136 808 25188 814
rect 25332 800 25360 1838
rect 25608 1358 25636 1838
rect 25596 1352 25648 1358
rect 25596 1294 25648 1300
rect 26068 882 26096 3878
rect 26252 2106 26280 4558
rect 26240 2100 26292 2106
rect 26240 2042 26292 2048
rect 26344 1986 26372 4626
rect 26516 4140 26568 4146
rect 26516 4082 26568 4088
rect 26424 3528 26476 3534
rect 26424 3470 26476 3476
rect 26252 1958 26372 1986
rect 26148 1896 26200 1902
rect 26148 1838 26200 1844
rect 26160 1494 26188 1838
rect 26148 1488 26200 1494
rect 26148 1430 26200 1436
rect 26056 876 26108 882
rect 26056 818 26108 824
rect 26252 800 26280 1958
rect 26436 1358 26464 3470
rect 26424 1352 26476 1358
rect 26424 1294 26476 1300
rect 26528 1018 26556 4082
rect 26608 3460 26660 3466
rect 26608 3402 26660 3408
rect 26620 2582 26648 3402
rect 26608 2576 26660 2582
rect 26608 2518 26660 2524
rect 26712 1358 26740 4966
rect 27344 4480 27396 4486
rect 27344 4422 27396 4428
rect 27356 3602 27384 4422
rect 27712 4072 27764 4078
rect 27712 4014 27764 4020
rect 27344 3596 27396 3602
rect 27344 3538 27396 3544
rect 26976 3392 27028 3398
rect 26976 3334 27028 3340
rect 27068 3392 27120 3398
rect 27068 3334 27120 3340
rect 26792 2372 26844 2378
rect 26792 2314 26844 2320
rect 26700 1352 26752 1358
rect 26700 1294 26752 1300
rect 26804 1170 26832 2314
rect 26988 1970 27016 3334
rect 27080 3194 27108 3334
rect 27068 3188 27120 3194
rect 27068 3130 27120 3136
rect 27620 3120 27672 3126
rect 27620 3062 27672 3068
rect 27160 2984 27212 2990
rect 27160 2926 27212 2932
rect 27068 2440 27120 2446
rect 27068 2382 27120 2388
rect 26884 1964 26936 1970
rect 26884 1906 26936 1912
rect 26976 1964 27028 1970
rect 26976 1906 27028 1912
rect 26896 1222 26924 1906
rect 26712 1142 26832 1170
rect 26884 1216 26936 1222
rect 26884 1158 26936 1164
rect 27080 1170 27108 2382
rect 27172 1358 27200 2926
rect 27528 2848 27580 2854
rect 27528 2790 27580 2796
rect 27540 2378 27568 2790
rect 27528 2372 27580 2378
rect 27528 2314 27580 2320
rect 27632 2106 27660 3062
rect 27724 2650 27752 4014
rect 27908 3738 27936 4966
rect 28080 4616 28132 4622
rect 28080 4558 28132 4564
rect 27896 3732 27948 3738
rect 27896 3674 27948 3680
rect 27896 3596 27948 3602
rect 27896 3538 27948 3544
rect 27804 3528 27856 3534
rect 27804 3470 27856 3476
rect 27712 2644 27764 2650
rect 27712 2586 27764 2592
rect 27620 2100 27672 2106
rect 27620 2042 27672 2048
rect 27816 1834 27844 3470
rect 27908 2990 27936 3538
rect 27988 3528 28040 3534
rect 27988 3470 28040 3476
rect 27896 2984 27948 2990
rect 27896 2926 27948 2932
rect 28000 2650 28028 3470
rect 28092 2854 28120 4558
rect 28172 2916 28224 2922
rect 28172 2858 28224 2864
rect 28080 2848 28132 2854
rect 28080 2790 28132 2796
rect 27988 2644 28040 2650
rect 27988 2586 28040 2592
rect 27804 1828 27856 1834
rect 27804 1770 27856 1776
rect 28184 1578 28212 2858
rect 28264 2440 28316 2446
rect 28264 2382 28316 2388
rect 28276 1834 28304 2382
rect 28264 1828 28316 1834
rect 28264 1770 28316 1776
rect 28092 1550 28212 1578
rect 27160 1352 27212 1358
rect 27160 1294 27212 1300
rect 27080 1142 27200 1170
rect 26516 1012 26568 1018
rect 26516 954 26568 960
rect 26712 800 26740 1142
rect 27172 800 27200 1142
rect 28092 800 28120 1550
rect 25136 750 25188 756
rect 25318 0 25374 800
rect 25778 0 25834 800
rect 26238 0 26294 800
rect 26698 0 26754 800
rect 27158 0 27214 800
rect 27618 0 27674 800
rect 28078 0 28134 800
rect 28368 746 28396 5102
rect 28632 4616 28684 4622
rect 28632 4558 28684 4564
rect 28448 3936 28500 3942
rect 28448 3878 28500 3884
rect 28460 2446 28488 3878
rect 28448 2440 28500 2446
rect 28448 2382 28500 2388
rect 28644 2310 28672 4558
rect 28920 2378 28948 5646
rect 29368 5568 29420 5574
rect 29368 5510 29420 5516
rect 29380 5234 29408 5510
rect 29184 5228 29236 5234
rect 29184 5170 29236 5176
rect 29368 5228 29420 5234
rect 29368 5170 29420 5176
rect 29196 4146 29224 5170
rect 29564 4758 29592 5646
rect 29552 4752 29604 4758
rect 29552 4694 29604 4700
rect 29276 4480 29328 4486
rect 29276 4422 29328 4428
rect 29288 4146 29316 4422
rect 29184 4140 29236 4146
rect 29184 4082 29236 4088
rect 29276 4140 29328 4146
rect 29276 4082 29328 4088
rect 29368 4072 29420 4078
rect 29368 4014 29420 4020
rect 29000 3936 29052 3942
rect 29000 3878 29052 3884
rect 29092 3936 29144 3942
rect 29092 3878 29144 3884
rect 28908 2372 28960 2378
rect 28908 2314 28960 2320
rect 28632 2304 28684 2310
rect 28632 2246 28684 2252
rect 29012 1970 29040 3878
rect 29104 3602 29132 3878
rect 29092 3596 29144 3602
rect 29092 3538 29144 3544
rect 29184 3392 29236 3398
rect 29184 3334 29236 3340
rect 29196 3126 29224 3334
rect 29184 3120 29236 3126
rect 29184 3062 29236 3068
rect 29276 2984 29328 2990
rect 29276 2926 29328 2932
rect 29000 1964 29052 1970
rect 29000 1906 29052 1912
rect 29288 1476 29316 2926
rect 29380 2650 29408 4014
rect 29564 2650 29592 4694
rect 29828 4616 29880 4622
rect 29828 4558 29880 4564
rect 29644 4548 29696 4554
rect 29644 4490 29696 4496
rect 29656 4146 29684 4490
rect 29644 4140 29696 4146
rect 29644 4082 29696 4088
rect 29840 3738 29868 4558
rect 30392 4078 30420 5646
rect 30656 5024 30708 5030
rect 30656 4966 30708 4972
rect 30472 4480 30524 4486
rect 30472 4422 30524 4428
rect 30564 4480 30616 4486
rect 30564 4422 30616 4428
rect 30484 4146 30512 4422
rect 30472 4140 30524 4146
rect 30472 4082 30524 4088
rect 30380 4072 30432 4078
rect 30380 4014 30432 4020
rect 29828 3732 29880 3738
rect 29828 3674 29880 3680
rect 29920 3732 29972 3738
rect 29920 3674 29972 3680
rect 29736 3664 29788 3670
rect 29736 3606 29788 3612
rect 29748 3516 29776 3606
rect 29748 3488 29868 3516
rect 29840 3058 29868 3488
rect 29828 3052 29880 3058
rect 29828 2994 29880 3000
rect 29368 2644 29420 2650
rect 29368 2586 29420 2592
rect 29552 2644 29604 2650
rect 29552 2586 29604 2592
rect 29288 1448 29500 1476
rect 29276 1352 29328 1358
rect 29276 1294 29328 1300
rect 28540 1284 28592 1290
rect 28540 1226 28592 1232
rect 28552 800 28580 1226
rect 29000 944 29052 950
rect 29000 886 29052 892
rect 29012 800 29040 886
rect 29288 814 29316 1294
rect 29276 808 29328 814
rect 28356 740 28408 746
rect 28356 682 28408 688
rect 28538 0 28594 800
rect 28998 0 29054 800
rect 29472 800 29500 1448
rect 29932 800 29960 3674
rect 30576 3466 30604 4422
rect 30668 4146 30696 4966
rect 30656 4140 30708 4146
rect 30656 4082 30708 4088
rect 30760 3738 30788 5646
rect 30840 5568 30892 5574
rect 30840 5510 30892 5516
rect 30748 3732 30800 3738
rect 30748 3674 30800 3680
rect 30564 3460 30616 3466
rect 30564 3402 30616 3408
rect 30748 3460 30800 3466
rect 30748 3402 30800 3408
rect 30104 3392 30156 3398
rect 30104 3334 30156 3340
rect 30012 2848 30064 2854
rect 30012 2790 30064 2796
rect 30024 2582 30052 2790
rect 30012 2576 30064 2582
rect 30012 2518 30064 2524
rect 30116 2514 30144 3334
rect 30472 2984 30524 2990
rect 30472 2926 30524 2932
rect 30484 2650 30512 2926
rect 30472 2644 30524 2650
rect 30472 2586 30524 2592
rect 30760 2514 30788 3402
rect 30104 2508 30156 2514
rect 30104 2450 30156 2456
rect 30748 2508 30800 2514
rect 30748 2450 30800 2456
rect 30380 1896 30432 1902
rect 30380 1838 30432 1844
rect 30392 800 30420 1838
rect 30852 1578 30880 5510
rect 31300 5160 31352 5166
rect 31300 5102 31352 5108
rect 31312 4826 31340 5102
rect 31300 4820 31352 4826
rect 31300 4762 31352 4768
rect 31300 4616 31352 4622
rect 31300 4558 31352 4564
rect 30932 4548 30984 4554
rect 30932 4490 30984 4496
rect 30944 3942 30972 4490
rect 31116 4208 31168 4214
rect 31116 4150 31168 4156
rect 31024 4072 31076 4078
rect 31024 4014 31076 4020
rect 30932 3936 30984 3942
rect 30932 3878 30984 3884
rect 31036 2446 31064 4014
rect 31128 2514 31156 4150
rect 31208 3936 31260 3942
rect 31208 3878 31260 3884
rect 31220 3058 31248 3878
rect 31208 3052 31260 3058
rect 31208 2994 31260 3000
rect 31116 2508 31168 2514
rect 31116 2450 31168 2456
rect 31024 2440 31076 2446
rect 31024 2382 31076 2388
rect 30760 1550 30880 1578
rect 30760 1290 30788 1550
rect 30840 1488 30892 1494
rect 30840 1430 30892 1436
rect 30748 1284 30800 1290
rect 30748 1226 30800 1232
rect 30472 1216 30524 1222
rect 30472 1158 30524 1164
rect 30484 1018 30512 1158
rect 30472 1012 30524 1018
rect 30472 954 30524 960
rect 30852 800 30880 1430
rect 31312 800 31340 4558
rect 31404 1766 31432 5646
rect 31576 5024 31628 5030
rect 31576 4966 31628 4972
rect 31392 1760 31444 1766
rect 31392 1702 31444 1708
rect 31588 1358 31616 4966
rect 31836 4922 32188 5972
rect 32312 5772 32364 5778
rect 32312 5714 32364 5720
rect 32220 5228 32272 5234
rect 32220 5170 32272 5176
rect 31836 4870 31858 4922
rect 31910 4870 31922 4922
rect 31974 4870 31986 4922
rect 32038 4870 32050 4922
rect 32102 4870 32114 4922
rect 32166 4870 32188 4922
rect 31836 3834 32188 4870
rect 31836 3782 31858 3834
rect 31910 3782 31922 3834
rect 31974 3782 31986 3834
rect 32038 3782 32050 3834
rect 32102 3782 32114 3834
rect 32166 3782 32188 3834
rect 31680 3454 31800 3482
rect 31680 3398 31708 3454
rect 31668 3392 31720 3398
rect 31668 3334 31720 3340
rect 31576 1352 31628 1358
rect 31576 1294 31628 1300
rect 31772 800 31800 3454
rect 31836 2746 32188 3782
rect 32232 3194 32260 5170
rect 32324 4146 32352 5714
rect 32864 5024 32916 5030
rect 32864 4966 32916 4972
rect 32680 4616 32732 4622
rect 32680 4558 32732 4564
rect 32404 4480 32456 4486
rect 32404 4422 32456 4428
rect 32312 4140 32364 4146
rect 32312 4082 32364 4088
rect 32312 3528 32364 3534
rect 32312 3470 32364 3476
rect 32220 3188 32272 3194
rect 32220 3130 32272 3136
rect 31836 2694 31858 2746
rect 31910 2694 31922 2746
rect 31974 2694 31986 2746
rect 32038 2694 32050 2746
rect 32102 2694 32114 2746
rect 32166 2694 32188 2746
rect 31836 2236 32188 2694
rect 32324 2650 32352 3470
rect 32312 2644 32364 2650
rect 32312 2586 32364 2592
rect 32416 2514 32444 4422
rect 32496 4072 32548 4078
rect 32496 4014 32548 4020
rect 32508 3194 32536 4014
rect 32588 3528 32640 3534
rect 32588 3470 32640 3476
rect 32600 3194 32628 3470
rect 32496 3188 32548 3194
rect 32496 3130 32548 3136
rect 32588 3188 32640 3194
rect 32588 3130 32640 3136
rect 32692 2582 32720 4558
rect 32876 4214 32904 4966
rect 32864 4208 32916 4214
rect 32864 4150 32916 4156
rect 32864 3936 32916 3942
rect 32864 3878 32916 3884
rect 32876 3602 32904 3878
rect 32864 3596 32916 3602
rect 32864 3538 32916 3544
rect 33060 3482 33088 7550
rect 36728 6520 36780 6526
rect 36728 6462 36780 6468
rect 34188 5466 34540 5972
rect 36740 5710 36768 6462
rect 42248 6316 42300 6322
rect 42248 6258 42300 6264
rect 41694 6080 41750 6089
rect 41694 6015 41750 6024
rect 39486 5944 39542 5953
rect 41708 5914 41736 6015
rect 39486 5879 39488 5888
rect 39540 5879 39542 5888
rect 41696 5908 41748 5914
rect 39488 5850 39540 5856
rect 41696 5850 41748 5856
rect 40408 5840 40460 5846
rect 40406 5808 40408 5817
rect 41604 5840 41656 5846
rect 40460 5808 40462 5817
rect 41604 5782 41656 5788
rect 40406 5743 40462 5752
rect 35164 5704 35216 5710
rect 35164 5646 35216 5652
rect 36452 5704 36504 5710
rect 36452 5646 36504 5652
rect 36728 5704 36780 5710
rect 36728 5646 36780 5652
rect 37188 5704 37240 5710
rect 37188 5646 37240 5652
rect 38108 5704 38160 5710
rect 38752 5704 38804 5710
rect 38108 5646 38160 5652
rect 38750 5672 38752 5681
rect 38844 5704 38896 5710
rect 38804 5672 38806 5681
rect 34188 5414 34210 5466
rect 34262 5414 34274 5466
rect 34326 5414 34338 5466
rect 34390 5414 34402 5466
rect 34454 5414 34466 5466
rect 34518 5414 34540 5466
rect 33416 5160 33468 5166
rect 33416 5102 33468 5108
rect 33784 5160 33836 5166
rect 33784 5102 33836 5108
rect 33140 4616 33192 4622
rect 33140 4558 33192 4564
rect 33152 4146 33180 4558
rect 33140 4140 33192 4146
rect 33140 4082 33192 4088
rect 33324 4140 33376 4146
rect 33324 4082 33376 4088
rect 33232 3936 33284 3942
rect 33232 3878 33284 3884
rect 32876 3454 33088 3482
rect 33140 3460 33192 3466
rect 32772 3392 32824 3398
rect 32772 3334 32824 3340
rect 32680 2576 32732 2582
rect 32680 2518 32732 2524
rect 32404 2508 32456 2514
rect 32404 2450 32456 2456
rect 31836 2180 31864 2236
rect 31920 2180 31944 2236
rect 32000 2180 32024 2236
rect 32080 2180 32104 2236
rect 32160 2180 32188 2236
rect 31836 2156 32188 2180
rect 31836 2100 31864 2156
rect 31920 2100 31944 2156
rect 32000 2100 32024 2156
rect 32080 2100 32104 2156
rect 32160 2100 32188 2156
rect 31836 2076 32188 2100
rect 31836 2020 31864 2076
rect 31920 2020 31944 2076
rect 32000 2020 32024 2076
rect 32080 2020 32104 2076
rect 32160 2020 32188 2076
rect 31836 1996 32188 2020
rect 31836 1940 31864 1996
rect 31920 1940 31944 1996
rect 32000 1940 32024 1996
rect 32080 1940 32104 1996
rect 32160 1940 32188 1996
rect 31836 1658 32188 1940
rect 32220 1896 32272 1902
rect 32784 1850 32812 3334
rect 32876 1970 32904 3454
rect 33140 3402 33192 3408
rect 32956 3392 33008 3398
rect 32956 3334 33008 3340
rect 33048 3392 33100 3398
rect 33048 3334 33100 3340
rect 32864 1964 32916 1970
rect 32864 1906 32916 1912
rect 32220 1838 32272 1844
rect 31836 1606 31858 1658
rect 31910 1606 31922 1658
rect 31974 1606 31986 1658
rect 32038 1606 32050 1658
rect 32102 1606 32114 1658
rect 32166 1606 32188 1658
rect 31836 1040 32188 1606
rect 32232 800 32260 1838
rect 32692 1822 32812 1850
rect 32692 800 32720 1822
rect 32968 1358 32996 3334
rect 33060 3058 33088 3334
rect 33048 3052 33100 3058
rect 33048 2994 33100 3000
rect 33048 2440 33100 2446
rect 33048 2382 33100 2388
rect 33060 1562 33088 2382
rect 33048 1556 33100 1562
rect 33048 1498 33100 1504
rect 32956 1352 33008 1358
rect 32956 1294 33008 1300
rect 33152 800 33180 3402
rect 33244 3058 33272 3878
rect 33232 3052 33284 3058
rect 33232 2994 33284 3000
rect 33336 2106 33364 4082
rect 33428 3738 33456 5102
rect 33796 4826 33824 5102
rect 33784 4820 33836 4826
rect 33784 4762 33836 4768
rect 33968 4616 34020 4622
rect 33968 4558 34020 4564
rect 34188 4588 34540 5414
rect 33876 4072 33928 4078
rect 33876 4014 33928 4020
rect 33416 3732 33468 3738
rect 33416 3674 33468 3680
rect 33692 3392 33744 3398
rect 33692 3334 33744 3340
rect 33784 3392 33836 3398
rect 33784 3334 33836 3340
rect 33704 3058 33732 3334
rect 33692 3052 33744 3058
rect 33692 2994 33744 3000
rect 33796 2514 33824 3334
rect 33784 2508 33836 2514
rect 33784 2450 33836 2456
rect 33324 2100 33376 2106
rect 33324 2042 33376 2048
rect 33508 1216 33560 1222
rect 33508 1158 33560 1164
rect 33520 864 33548 1158
rect 33888 1018 33916 4014
rect 33980 2854 34008 4558
rect 34188 4532 34216 4588
rect 34272 4532 34296 4588
rect 34352 4532 34376 4588
rect 34432 4532 34456 4588
rect 34512 4532 34540 4588
rect 34612 4616 34664 4622
rect 34612 4558 34664 4564
rect 34188 4508 34540 4532
rect 34188 4452 34216 4508
rect 34272 4452 34296 4508
rect 34352 4452 34376 4508
rect 34432 4452 34456 4508
rect 34512 4452 34540 4508
rect 34188 4428 34540 4452
rect 34188 4378 34216 4428
rect 34272 4378 34296 4428
rect 34352 4378 34376 4428
rect 34432 4378 34456 4428
rect 34512 4378 34540 4428
rect 34188 4326 34210 4378
rect 34272 4372 34274 4378
rect 34454 4372 34456 4378
rect 34262 4348 34274 4372
rect 34326 4348 34338 4372
rect 34390 4348 34402 4372
rect 34454 4348 34466 4372
rect 34272 4326 34274 4348
rect 34454 4326 34456 4348
rect 34518 4326 34540 4378
rect 34188 4292 34216 4326
rect 34272 4292 34296 4326
rect 34352 4292 34376 4326
rect 34432 4292 34456 4326
rect 34512 4292 34540 4326
rect 34060 3936 34112 3942
rect 34060 3878 34112 3884
rect 34072 3602 34100 3878
rect 34060 3596 34112 3602
rect 34060 3538 34112 3544
rect 34188 3290 34540 4292
rect 34188 3238 34210 3290
rect 34262 3238 34274 3290
rect 34326 3238 34338 3290
rect 34390 3238 34402 3290
rect 34454 3238 34466 3290
rect 34518 3238 34540 3290
rect 33968 2848 34020 2854
rect 33968 2790 34020 2796
rect 34188 2202 34540 3238
rect 34624 2650 34652 4558
rect 34796 4072 34848 4078
rect 34796 4014 34848 4020
rect 34980 4072 35032 4078
rect 34980 4014 35032 4020
rect 34704 3528 34756 3534
rect 34704 3470 34756 3476
rect 34612 2644 34664 2650
rect 34612 2586 34664 2592
rect 34716 2582 34744 3470
rect 34808 2666 34836 4014
rect 34888 3392 34940 3398
rect 34888 3334 34940 3340
rect 34900 3058 34928 3334
rect 34992 3194 35020 4014
rect 35072 3936 35124 3942
rect 35072 3878 35124 3884
rect 34980 3188 35032 3194
rect 34980 3130 35032 3136
rect 34888 3052 34940 3058
rect 34888 2994 34940 3000
rect 34980 2984 35032 2990
rect 34980 2926 35032 2932
rect 34808 2638 34928 2666
rect 34704 2576 34756 2582
rect 34704 2518 34756 2524
rect 34796 2576 34848 2582
rect 34796 2518 34848 2524
rect 34612 2372 34664 2378
rect 34612 2314 34664 2320
rect 34188 2150 34210 2202
rect 34262 2150 34274 2202
rect 34326 2150 34338 2202
rect 34390 2150 34402 2202
rect 34454 2150 34466 2202
rect 34518 2150 34540 2202
rect 34060 1896 34112 1902
rect 34060 1838 34112 1844
rect 33968 1284 34020 1290
rect 33968 1226 34020 1232
rect 33876 1012 33928 1018
rect 33876 954 33928 960
rect 33980 950 34008 1226
rect 33968 944 34020 950
rect 33968 886 34020 892
rect 33520 836 33640 864
rect 33612 800 33640 836
rect 34072 800 34100 1838
rect 34188 1114 34540 2150
rect 34188 1062 34210 1114
rect 34262 1062 34274 1114
rect 34326 1062 34338 1114
rect 34390 1062 34402 1114
rect 34454 1062 34466 1114
rect 34518 1062 34540 1114
rect 34188 1040 34540 1062
rect 34624 898 34652 2314
rect 34808 1970 34836 2518
rect 34900 2310 34928 2638
rect 34888 2304 34940 2310
rect 34888 2246 34940 2252
rect 34796 1964 34848 1970
rect 34796 1906 34848 1912
rect 34532 870 34652 898
rect 34532 800 34560 870
rect 34992 800 35020 2926
rect 35084 1290 35112 3878
rect 35176 3466 35204 5646
rect 36464 5370 36492 5646
rect 36452 5364 36504 5370
rect 36452 5306 36504 5312
rect 36544 5160 36596 5166
rect 36544 5102 36596 5108
rect 36084 5024 36136 5030
rect 36084 4966 36136 4972
rect 36096 4690 36124 4966
rect 36084 4684 36136 4690
rect 36084 4626 36136 4632
rect 36360 4616 36412 4622
rect 36360 4558 36412 4564
rect 35256 4548 35308 4554
rect 35256 4490 35308 4496
rect 35268 3738 35296 4490
rect 35992 4072 36044 4078
rect 35992 4014 36044 4020
rect 35256 3732 35308 3738
rect 35256 3674 35308 3680
rect 35900 3528 35952 3534
rect 35900 3470 35952 3476
rect 35164 3460 35216 3466
rect 35164 3402 35216 3408
rect 35624 3460 35676 3466
rect 35624 3402 35676 3408
rect 35636 3058 35664 3402
rect 35624 3052 35676 3058
rect 35624 2994 35676 3000
rect 35532 2440 35584 2446
rect 35532 2382 35584 2388
rect 35544 1562 35572 2382
rect 35716 2304 35768 2310
rect 35716 2246 35768 2252
rect 35728 1970 35756 2246
rect 35624 1964 35676 1970
rect 35624 1906 35676 1912
rect 35716 1964 35768 1970
rect 35716 1906 35768 1912
rect 35532 1556 35584 1562
rect 35532 1498 35584 1504
rect 35636 1494 35664 1906
rect 35624 1488 35676 1494
rect 35624 1430 35676 1436
rect 35072 1284 35124 1290
rect 35072 1226 35124 1232
rect 35440 1284 35492 1290
rect 35440 1226 35492 1232
rect 35452 800 35480 1226
rect 35912 800 35940 3470
rect 36004 3194 36032 4014
rect 36084 3528 36136 3534
rect 36084 3470 36136 3476
rect 35992 3188 36044 3194
rect 35992 3130 36044 3136
rect 36096 2650 36124 3470
rect 36372 3194 36400 4558
rect 36360 3188 36412 3194
rect 36360 3130 36412 3136
rect 36176 2848 36228 2854
rect 36176 2790 36228 2796
rect 36084 2644 36136 2650
rect 36084 2586 36136 2592
rect 36188 2514 36216 2790
rect 36176 2508 36228 2514
rect 36176 2450 36228 2456
rect 36360 2440 36412 2446
rect 36360 2382 36412 2388
rect 36268 2372 36320 2378
rect 36268 2314 36320 2320
rect 36280 2106 36308 2314
rect 36268 2100 36320 2106
rect 36268 2042 36320 2048
rect 36372 800 36400 2382
rect 36556 2038 36584 5102
rect 36912 4548 36964 4554
rect 36912 4490 36964 4496
rect 36728 4480 36780 4486
rect 36728 4422 36780 4428
rect 36740 4282 36768 4422
rect 36728 4276 36780 4282
rect 36728 4218 36780 4224
rect 36820 3936 36872 3942
rect 36820 3878 36872 3884
rect 36832 3058 36860 3878
rect 36820 3052 36872 3058
rect 36820 2994 36872 3000
rect 36924 2650 36952 4490
rect 37200 4010 37228 5646
rect 37280 5568 37332 5574
rect 37280 5510 37332 5516
rect 37292 5234 37320 5510
rect 38120 5302 38148 5646
rect 38844 5646 38896 5652
rect 39764 5704 39816 5710
rect 39764 5646 39816 5652
rect 40408 5704 40460 5710
rect 40408 5646 40460 5652
rect 38750 5607 38806 5616
rect 38108 5296 38160 5302
rect 38108 5238 38160 5244
rect 37280 5228 37332 5234
rect 37280 5170 37332 5176
rect 37740 5160 37792 5166
rect 37740 5102 37792 5108
rect 37752 4622 37780 5102
rect 38856 5030 38884 5646
rect 38936 5636 38988 5642
rect 38936 5578 38988 5584
rect 38844 5024 38896 5030
rect 38844 4966 38896 4972
rect 37740 4616 37792 4622
rect 37740 4558 37792 4564
rect 38016 4548 38068 4554
rect 38016 4490 38068 4496
rect 37924 4480 37976 4486
rect 37924 4422 37976 4428
rect 37936 4214 37964 4422
rect 37924 4208 37976 4214
rect 37924 4150 37976 4156
rect 37832 4140 37884 4146
rect 37832 4082 37884 4088
rect 37188 4004 37240 4010
rect 37188 3946 37240 3952
rect 37464 3392 37516 3398
rect 37464 3334 37516 3340
rect 37280 2984 37332 2990
rect 37280 2926 37332 2932
rect 36912 2644 36964 2650
rect 36912 2586 36964 2592
rect 37292 2106 37320 2926
rect 37280 2100 37332 2106
rect 37280 2042 37332 2048
rect 36544 2032 36596 2038
rect 36544 1974 36596 1980
rect 37476 1970 37504 3334
rect 37844 2514 37872 4082
rect 38028 3194 38056 4490
rect 38948 4146 38976 5578
rect 39212 5160 39264 5166
rect 39210 5128 39212 5137
rect 39264 5128 39266 5137
rect 39210 5063 39266 5072
rect 38936 4140 38988 4146
rect 38936 4082 38988 4088
rect 38384 3528 38436 3534
rect 38384 3470 38436 3476
rect 39120 3528 39172 3534
rect 39120 3470 39172 3476
rect 38016 3188 38068 3194
rect 38016 3130 38068 3136
rect 38396 2650 38424 3470
rect 38752 2848 38804 2854
rect 38752 2790 38804 2796
rect 38384 2644 38436 2650
rect 38384 2586 38436 2592
rect 38764 2514 38792 2790
rect 37832 2508 37884 2514
rect 37832 2450 37884 2456
rect 38752 2508 38804 2514
rect 38752 2450 38804 2456
rect 37648 2440 37700 2446
rect 37700 2400 37780 2428
rect 37648 2382 37700 2388
rect 37464 1964 37516 1970
rect 37464 1906 37516 1912
rect 36820 1896 36872 1902
rect 36820 1838 36872 1844
rect 36544 1284 36596 1290
rect 36544 1226 36596 1232
rect 36556 1018 36584 1226
rect 36544 1012 36596 1018
rect 36544 954 36596 960
rect 36832 800 36860 1838
rect 36912 1352 36964 1358
rect 36912 1294 36964 1300
rect 29276 750 29328 756
rect 29458 0 29514 800
rect 29918 0 29974 800
rect 30378 0 30434 800
rect 30838 0 30894 800
rect 31298 0 31354 800
rect 31758 0 31814 800
rect 32218 0 32274 800
rect 32678 0 32734 800
rect 33138 0 33194 800
rect 33598 0 33654 800
rect 34058 0 34114 800
rect 34518 0 34574 800
rect 34978 0 35034 800
rect 35438 0 35494 800
rect 35898 0 35954 800
rect 36358 0 36414 800
rect 36818 0 36874 800
rect 36924 678 36952 1294
rect 37280 1284 37332 1290
rect 37280 1226 37332 1232
rect 37292 800 37320 1226
rect 37752 800 37780 2400
rect 39132 2106 39160 3470
rect 39580 2304 39632 2310
rect 39580 2246 39632 2252
rect 39120 2100 39172 2106
rect 39120 2042 39172 2048
rect 39592 1970 39620 2246
rect 39580 1964 39632 1970
rect 39580 1906 39632 1912
rect 39120 1896 39172 1902
rect 39120 1838 39172 1844
rect 38660 1420 38712 1426
rect 38660 1362 38712 1368
rect 38200 1284 38252 1290
rect 38200 1226 38252 1232
rect 38212 800 38240 1226
rect 38672 800 38700 1362
rect 39132 800 39160 1838
rect 39396 1352 39448 1358
rect 39396 1294 39448 1300
rect 36912 672 36964 678
rect 36912 614 36964 620
rect 37278 0 37334 800
rect 37738 0 37794 800
rect 38198 0 38254 800
rect 38658 0 38714 800
rect 39118 0 39174 800
rect 39408 610 39436 1294
rect 39580 1284 39632 1290
rect 39580 1226 39632 1232
rect 39592 800 39620 1226
rect 39776 1018 39804 5646
rect 40132 5160 40184 5166
rect 40132 5102 40184 5108
rect 39948 5092 40000 5098
rect 39948 5034 40000 5040
rect 39960 4622 39988 5034
rect 39948 4616 40000 4622
rect 39948 4558 40000 4564
rect 40144 3738 40172 5102
rect 40224 4616 40276 4622
rect 40224 4558 40276 4564
rect 40132 3732 40184 3738
rect 40132 3674 40184 3680
rect 40236 3126 40264 4558
rect 40314 3632 40370 3641
rect 40314 3567 40370 3576
rect 40328 3534 40356 3567
rect 40316 3528 40368 3534
rect 40316 3470 40368 3476
rect 40224 3120 40276 3126
rect 40224 3062 40276 3068
rect 39856 3052 39908 3058
rect 39856 2994 39908 3000
rect 40040 3052 40092 3058
rect 40040 2994 40092 3000
rect 39868 2106 39896 2994
rect 39856 2100 39908 2106
rect 39856 2042 39908 2048
rect 39764 1012 39816 1018
rect 39764 954 39816 960
rect 40052 800 40080 2994
rect 40132 2984 40184 2990
rect 40132 2926 40184 2932
rect 40224 2984 40276 2990
rect 40224 2926 40276 2932
rect 40144 1290 40172 2926
rect 40236 2650 40264 2926
rect 40224 2644 40276 2650
rect 40224 2586 40276 2592
rect 40316 2304 40368 2310
rect 40316 2246 40368 2252
rect 40328 1970 40356 2246
rect 40316 1964 40368 1970
rect 40316 1906 40368 1912
rect 40132 1284 40184 1290
rect 40132 1226 40184 1232
rect 40420 950 40448 5646
rect 41616 5370 41644 5782
rect 41604 5364 41656 5370
rect 41604 5306 41656 5312
rect 41836 4922 42188 5972
rect 42260 5302 42288 6258
rect 42708 5704 42760 5710
rect 42708 5646 42760 5652
rect 42720 5370 42748 5646
rect 44188 5466 44540 5972
rect 44732 5772 44784 5778
rect 44732 5714 44784 5720
rect 44188 5414 44210 5466
rect 44262 5414 44274 5466
rect 44326 5414 44338 5466
rect 44390 5414 44402 5466
rect 44454 5414 44466 5466
rect 44518 5414 44540 5466
rect 42708 5364 42760 5370
rect 42708 5306 42760 5312
rect 42892 5364 42944 5370
rect 42892 5306 42944 5312
rect 42248 5296 42300 5302
rect 42248 5238 42300 5244
rect 41836 4870 41858 4922
rect 41910 4870 41922 4922
rect 41974 4870 41986 4922
rect 42038 4870 42050 4922
rect 42102 4870 42114 4922
rect 42166 4870 42188 4922
rect 40590 4856 40646 4865
rect 40590 4791 40646 4800
rect 40604 4758 40632 4791
rect 40592 4752 40644 4758
rect 40592 4694 40644 4700
rect 41326 4040 41382 4049
rect 41326 3975 41328 3984
rect 41380 3975 41382 3984
rect 41328 3946 41380 3952
rect 41512 3936 41564 3942
rect 41512 3878 41564 3884
rect 40866 3768 40922 3777
rect 40866 3703 40922 3712
rect 40880 3670 40908 3703
rect 40868 3664 40920 3670
rect 40868 3606 40920 3612
rect 41524 3602 41552 3878
rect 41836 3834 42188 4870
rect 42248 4072 42300 4078
rect 42248 4014 42300 4020
rect 41836 3782 41858 3834
rect 41910 3782 41922 3834
rect 41974 3782 41986 3834
rect 42038 3782 42050 3834
rect 42102 3782 42114 3834
rect 42166 3782 42188 3834
rect 41512 3596 41564 3602
rect 41512 3538 41564 3544
rect 40592 3528 40644 3534
rect 40592 3470 40644 3476
rect 41328 3528 41380 3534
rect 41328 3470 41380 3476
rect 41604 3528 41656 3534
rect 41604 3470 41656 3476
rect 40604 2106 40632 3470
rect 41052 2440 41104 2446
rect 41052 2382 41104 2388
rect 40776 2372 40828 2378
rect 40776 2314 40828 2320
rect 40592 2100 40644 2106
rect 40592 2042 40644 2048
rect 40500 1760 40552 1766
rect 40500 1702 40552 1708
rect 40512 1358 40540 1702
rect 40500 1352 40552 1358
rect 40500 1294 40552 1300
rect 40408 944 40460 950
rect 40408 886 40460 892
rect 40512 870 40632 898
rect 40512 800 40540 870
rect 39396 604 39448 610
rect 39396 546 39448 552
rect 39578 0 39634 800
rect 40038 0 40094 800
rect 40498 0 40554 800
rect 40604 762 40632 870
rect 40788 762 40816 2314
rect 41064 1222 41092 2382
rect 41340 1562 41368 3470
rect 41420 2848 41472 2854
rect 41420 2790 41472 2796
rect 41512 2848 41564 2854
rect 41512 2790 41564 2796
rect 41432 1970 41460 2790
rect 41524 2514 41552 2790
rect 41512 2508 41564 2514
rect 41512 2450 41564 2456
rect 41420 1964 41472 1970
rect 41420 1906 41472 1912
rect 41328 1556 41380 1562
rect 41328 1498 41380 1504
rect 41616 1442 41644 3470
rect 41694 2952 41750 2961
rect 41694 2887 41696 2896
rect 41748 2887 41750 2896
rect 41696 2858 41748 2864
rect 41432 1414 41644 1442
rect 41836 2746 42188 3782
rect 42260 3738 42288 4014
rect 42248 3732 42300 3738
rect 42248 3674 42300 3680
rect 42248 3596 42300 3602
rect 42248 3538 42300 3544
rect 41836 2694 41858 2746
rect 41910 2694 41922 2746
rect 41974 2694 41986 2746
rect 42038 2694 42050 2746
rect 42102 2694 42114 2746
rect 42166 2694 42188 2746
rect 41836 2236 42188 2694
rect 41836 2180 41864 2236
rect 41920 2180 41944 2236
rect 42000 2180 42024 2236
rect 42080 2180 42104 2236
rect 42160 2180 42188 2236
rect 41836 2156 42188 2180
rect 41836 2100 41864 2156
rect 41920 2100 41944 2156
rect 42000 2100 42024 2156
rect 42080 2100 42104 2156
rect 42160 2100 42188 2156
rect 41836 2076 42188 2100
rect 41836 2020 41864 2076
rect 41920 2020 41944 2076
rect 42000 2020 42024 2076
rect 42080 2020 42104 2076
rect 42160 2020 42188 2076
rect 41836 1996 42188 2020
rect 41836 1940 41864 1996
rect 41920 1940 41944 1996
rect 42000 1940 42024 1996
rect 42080 1940 42104 1996
rect 42160 1940 42188 1996
rect 41836 1658 42188 1940
rect 41836 1606 41858 1658
rect 41910 1606 41922 1658
rect 41974 1606 41986 1658
rect 42038 1606 42050 1658
rect 42102 1606 42114 1658
rect 42166 1606 42188 1658
rect 41144 1352 41196 1358
rect 41144 1294 41196 1300
rect 41052 1216 41104 1222
rect 41052 1158 41104 1164
rect 41156 1018 41184 1294
rect 41328 1284 41380 1290
rect 41328 1226 41380 1232
rect 41144 1012 41196 1018
rect 41144 954 41196 960
rect 40972 870 41092 898
rect 40972 800 41000 870
rect 40604 734 40816 762
rect 40958 0 41014 800
rect 41064 762 41092 870
rect 41340 762 41368 1226
rect 41432 800 41460 1414
rect 41836 1040 42188 1606
rect 41892 870 42012 898
rect 41892 800 41920 870
rect 41064 734 41368 762
rect 41418 0 41474 800
rect 41878 0 41934 800
rect 41984 762 42012 870
rect 42260 762 42288 3538
rect 42340 3460 42392 3466
rect 42340 3402 42392 3408
rect 42352 3194 42380 3402
rect 42524 3392 42576 3398
rect 42524 3334 42576 3340
rect 42340 3188 42392 3194
rect 42340 3130 42392 3136
rect 42338 3088 42394 3097
rect 42338 3023 42394 3032
rect 42352 2854 42380 3023
rect 42340 2848 42392 2854
rect 42340 2790 42392 2796
rect 42536 2514 42564 3334
rect 42720 2961 42748 5306
rect 42904 4486 42932 5306
rect 44086 5264 44142 5273
rect 44086 5199 44088 5208
rect 44140 5199 44142 5208
rect 44088 5170 44140 5176
rect 43628 5092 43680 5098
rect 43628 5034 43680 5040
rect 43640 4758 43668 5034
rect 43628 4752 43680 4758
rect 43628 4694 43680 4700
rect 44088 4616 44140 4622
rect 44088 4558 44140 4564
rect 44188 4588 44540 5414
rect 44744 5234 44772 5714
rect 44732 5228 44784 5234
rect 44732 5170 44784 5176
rect 44836 4622 44864 7686
rect 46756 6384 46808 6390
rect 46756 6326 46808 6332
rect 45468 5568 45520 5574
rect 45468 5510 45520 5516
rect 45480 5234 45508 5510
rect 46112 5296 46164 5302
rect 46112 5238 46164 5244
rect 46202 5264 46258 5273
rect 45468 5228 45520 5234
rect 45468 5170 45520 5176
rect 42892 4480 42944 4486
rect 42892 4422 42944 4428
rect 43536 4276 43588 4282
rect 43536 4218 43588 4224
rect 43548 4146 43576 4218
rect 43536 4140 43588 4146
rect 43536 4082 43588 4088
rect 43352 4072 43404 4078
rect 44100 4049 44128 4558
rect 44188 4532 44216 4588
rect 44272 4532 44296 4588
rect 44352 4532 44376 4588
rect 44432 4532 44456 4588
rect 44512 4532 44540 4588
rect 44824 4616 44876 4622
rect 44824 4558 44876 4564
rect 45008 4616 45060 4622
rect 45008 4558 45060 4564
rect 45100 4616 45152 4622
rect 45100 4558 45152 4564
rect 44188 4508 44540 4532
rect 44188 4452 44216 4508
rect 44272 4452 44296 4508
rect 44352 4452 44376 4508
rect 44432 4452 44456 4508
rect 44512 4452 44540 4508
rect 44188 4428 44540 4452
rect 44188 4378 44216 4428
rect 44272 4378 44296 4428
rect 44352 4378 44376 4428
rect 44432 4378 44456 4428
rect 44512 4378 44540 4428
rect 44188 4326 44210 4378
rect 44272 4372 44274 4378
rect 44454 4372 44456 4378
rect 44262 4348 44274 4372
rect 44326 4348 44338 4372
rect 44390 4348 44402 4372
rect 44454 4348 44466 4372
rect 44272 4326 44274 4348
rect 44454 4326 44456 4348
rect 44518 4326 44540 4378
rect 44188 4292 44216 4326
rect 44272 4292 44296 4326
rect 44352 4292 44376 4326
rect 44432 4292 44456 4326
rect 44512 4292 44540 4326
rect 43352 4014 43404 4020
rect 44086 4040 44142 4049
rect 43364 3738 43392 4014
rect 44086 3975 44142 3984
rect 43812 3936 43864 3942
rect 43812 3878 43864 3884
rect 43352 3732 43404 3738
rect 43352 3674 43404 3680
rect 43444 3392 43496 3398
rect 43444 3334 43496 3340
rect 43536 3392 43588 3398
rect 43536 3334 43588 3340
rect 42984 2984 43036 2990
rect 42706 2952 42762 2961
rect 42984 2926 43036 2932
rect 42706 2887 42762 2896
rect 42996 2650 43024 2926
rect 42984 2644 43036 2650
rect 42984 2586 43036 2592
rect 43456 2514 43484 3334
rect 43548 3126 43576 3334
rect 43536 3120 43588 3126
rect 43536 3062 43588 3068
rect 43824 3058 43852 3878
rect 44188 3290 44540 4292
rect 45020 3670 45048 4558
rect 45008 3664 45060 3670
rect 45112 3641 45140 4558
rect 45652 4480 45704 4486
rect 45652 4422 45704 4428
rect 45664 4282 45692 4422
rect 45652 4276 45704 4282
rect 45652 4218 45704 4224
rect 46124 4214 46152 5238
rect 46202 5199 46204 5208
rect 46256 5199 46258 5208
rect 46204 5170 46256 5176
rect 46664 5160 46716 5166
rect 46662 5128 46664 5137
rect 46716 5128 46718 5137
rect 46662 5063 46718 5072
rect 46768 4622 46796 6326
rect 47320 5370 47348 7754
rect 55784 7478 55812 7754
rect 55772 7472 55824 7478
rect 55772 7414 55824 7420
rect 63132 7472 63184 7478
rect 63132 7414 63184 7420
rect 62672 7404 62724 7410
rect 62672 7346 62724 7352
rect 62304 7336 62356 7342
rect 62304 7278 62356 7284
rect 55036 7268 55088 7274
rect 55036 7210 55088 7216
rect 49056 6860 49108 6866
rect 49056 6802 49108 6808
rect 47768 6656 47820 6662
rect 47768 6598 47820 6604
rect 47308 5364 47360 5370
rect 47308 5306 47360 5312
rect 47584 5160 47636 5166
rect 47584 5102 47636 5108
rect 47596 4865 47624 5102
rect 47582 4856 47638 4865
rect 47582 4791 47638 4800
rect 47780 4622 47808 6598
rect 48228 6452 48280 6458
rect 48228 6394 48280 6400
rect 48240 5370 48268 6394
rect 48964 5704 49016 5710
rect 48964 5646 49016 5652
rect 48228 5364 48280 5370
rect 48228 5306 48280 5312
rect 48976 5302 49004 5646
rect 49068 5370 49096 6802
rect 49792 6792 49844 6798
rect 49792 6734 49844 6740
rect 49608 6588 49660 6594
rect 49608 6530 49660 6536
rect 49620 5914 49648 6530
rect 49608 5908 49660 5914
rect 49608 5850 49660 5856
rect 49700 5704 49752 5710
rect 49700 5646 49752 5652
rect 49056 5364 49108 5370
rect 49056 5306 49108 5312
rect 48964 5296 49016 5302
rect 48964 5238 49016 5244
rect 48412 5160 48464 5166
rect 48412 5102 48464 5108
rect 49148 5160 49200 5166
rect 49148 5102 49200 5108
rect 46756 4616 46808 4622
rect 46756 4558 46808 4564
rect 47216 4616 47268 4622
rect 47216 4558 47268 4564
rect 47768 4616 47820 4622
rect 47768 4558 47820 4564
rect 47860 4616 47912 4622
rect 47860 4558 47912 4564
rect 46112 4208 46164 4214
rect 46112 4150 46164 4156
rect 45468 4072 45520 4078
rect 45468 4014 45520 4020
rect 45008 3606 45060 3612
rect 45098 3632 45154 3641
rect 44732 3596 44784 3602
rect 45098 3567 45154 3576
rect 44732 3538 44784 3544
rect 44640 3528 44692 3534
rect 44640 3470 44692 3476
rect 44188 3238 44210 3290
rect 44262 3238 44274 3290
rect 44326 3238 44338 3290
rect 44390 3238 44402 3290
rect 44454 3238 44466 3290
rect 44518 3238 44540 3290
rect 43812 3052 43864 3058
rect 43812 2994 43864 3000
rect 42524 2508 42576 2514
rect 42524 2450 42576 2456
rect 43444 2508 43496 2514
rect 43444 2450 43496 2456
rect 44188 2202 44540 3238
rect 44652 3194 44680 3470
rect 44640 3188 44692 3194
rect 44640 3130 44692 3136
rect 44640 2984 44692 2990
rect 44640 2926 44692 2932
rect 44652 2650 44680 2926
rect 44640 2644 44692 2650
rect 44640 2586 44692 2592
rect 44188 2150 44210 2202
rect 44262 2150 44274 2202
rect 44326 2150 44338 2202
rect 44390 2150 44402 2202
rect 44454 2150 44466 2202
rect 44518 2150 44540 2202
rect 42340 1896 42392 1902
rect 42340 1838 42392 1844
rect 43720 1896 43772 1902
rect 43720 1838 43772 1844
rect 42352 800 42380 1838
rect 43260 1760 43312 1766
rect 43260 1702 43312 1708
rect 42800 1420 42852 1426
rect 42800 1362 42852 1368
rect 42812 800 42840 1362
rect 43272 800 43300 1702
rect 43732 800 43760 1838
rect 43996 1352 44048 1358
rect 43996 1294 44048 1300
rect 44008 882 44036 1294
rect 44188 1114 44540 2150
rect 44744 1442 44772 3538
rect 45480 3398 45508 4014
rect 45560 3528 45612 3534
rect 45560 3470 45612 3476
rect 45468 3392 45520 3398
rect 45468 3334 45520 3340
rect 45376 2916 45428 2922
rect 45376 2858 45428 2864
rect 44824 2304 44876 2310
rect 44824 2246 44876 2252
rect 44916 2304 44968 2310
rect 44916 2246 44968 2252
rect 44188 1062 44210 1114
rect 44262 1062 44274 1114
rect 44326 1062 44338 1114
rect 44390 1062 44402 1114
rect 44454 1062 44466 1114
rect 44518 1062 44540 1114
rect 44188 1040 44540 1062
rect 44652 1414 44772 1442
rect 43996 876 44048 882
rect 43996 818 44048 824
rect 44652 800 44680 1414
rect 44836 1358 44864 2246
rect 44928 1970 44956 2246
rect 45388 2106 45416 2858
rect 45572 2650 45600 3470
rect 47124 3460 47176 3466
rect 47124 3402 47176 3408
rect 46940 3392 46992 3398
rect 46940 3334 46992 3340
rect 47032 3392 47084 3398
rect 47032 3334 47084 3340
rect 46112 2984 46164 2990
rect 46112 2926 46164 2932
rect 46848 2984 46900 2990
rect 46848 2926 46900 2932
rect 46020 2916 46072 2922
rect 46020 2858 46072 2864
rect 45928 2848 45980 2854
rect 45928 2790 45980 2796
rect 45560 2644 45612 2650
rect 45560 2586 45612 2592
rect 45560 2440 45612 2446
rect 45560 2382 45612 2388
rect 45376 2100 45428 2106
rect 45376 2042 45428 2048
rect 44916 1964 44968 1970
rect 44916 1906 44968 1912
rect 45572 1562 45600 2382
rect 45940 1970 45968 2790
rect 45928 1964 45980 1970
rect 45928 1906 45980 1912
rect 45560 1556 45612 1562
rect 45560 1498 45612 1504
rect 44824 1352 44876 1358
rect 44824 1294 44876 1300
rect 45100 1284 45152 1290
rect 45100 1226 45152 1232
rect 45112 800 45140 1226
rect 46032 800 46060 2858
rect 46124 2650 46152 2926
rect 46112 2644 46164 2650
rect 46112 2586 46164 2592
rect 46112 2440 46164 2446
rect 46112 2382 46164 2388
rect 46124 2106 46152 2382
rect 46112 2100 46164 2106
rect 46112 2042 46164 2048
rect 46860 1970 46888 2926
rect 46952 2514 46980 3334
rect 46940 2508 46992 2514
rect 46940 2450 46992 2456
rect 46940 2304 46992 2310
rect 46940 2246 46992 2252
rect 46848 1964 46900 1970
rect 46848 1906 46900 1912
rect 46664 1896 46716 1902
rect 46664 1838 46716 1844
rect 46676 1766 46704 1838
rect 46664 1760 46716 1766
rect 46664 1702 46716 1708
rect 46952 1562 46980 2246
rect 47044 1970 47072 3334
rect 47136 2514 47164 3402
rect 47124 2508 47176 2514
rect 47124 2450 47176 2456
rect 47228 2378 47256 4558
rect 47584 4072 47636 4078
rect 47768 4072 47820 4078
rect 47636 4032 47768 4060
rect 47584 4014 47636 4020
rect 47768 4014 47820 4020
rect 47872 3777 47900 4558
rect 47952 4140 48004 4146
rect 47952 4082 48004 4088
rect 47858 3768 47914 3777
rect 47858 3703 47914 3712
rect 47492 3528 47544 3534
rect 47492 3470 47544 3476
rect 47504 3194 47532 3470
rect 47492 3188 47544 3194
rect 47492 3130 47544 3136
rect 47964 3097 47992 4082
rect 48424 3738 48452 5102
rect 49160 4826 49188 5102
rect 49148 4820 49200 4826
rect 49148 4762 49200 4768
rect 49712 4706 49740 5646
rect 49804 5370 49832 6734
rect 50712 6248 50764 6254
rect 50712 6190 50764 6196
rect 50724 5914 50752 6190
rect 50712 5908 50764 5914
rect 50712 5850 50764 5856
rect 50804 5704 50856 5710
rect 50804 5646 50856 5652
rect 51540 5704 51592 5710
rect 51540 5646 51592 5652
rect 49792 5364 49844 5370
rect 49792 5306 49844 5312
rect 49792 5160 49844 5166
rect 49792 5102 49844 5108
rect 50160 5160 50212 5166
rect 50160 5102 50212 5108
rect 49344 4678 49740 4706
rect 49344 4078 49372 4678
rect 49608 4616 49660 4622
rect 49608 4558 49660 4564
rect 49332 4072 49384 4078
rect 49332 4014 49384 4020
rect 49424 4072 49476 4078
rect 49424 4014 49476 4020
rect 49436 3738 49464 4014
rect 49620 3890 49648 4558
rect 49528 3862 49648 3890
rect 48412 3732 48464 3738
rect 48412 3674 48464 3680
rect 49424 3732 49476 3738
rect 49424 3674 49476 3680
rect 48320 3664 48372 3670
rect 48320 3606 48372 3612
rect 47950 3088 48006 3097
rect 47950 3023 48006 3032
rect 47400 2848 47452 2854
rect 47400 2790 47452 2796
rect 47308 2508 47360 2514
rect 47308 2450 47360 2456
rect 47216 2372 47268 2378
rect 47216 2314 47268 2320
rect 47032 1964 47084 1970
rect 47032 1906 47084 1912
rect 47320 1766 47348 2450
rect 47308 1760 47360 1766
rect 47308 1702 47360 1708
rect 46940 1556 46992 1562
rect 46940 1498 46992 1504
rect 46388 1352 46440 1358
rect 46388 1294 46440 1300
rect 41984 734 42288 762
rect 42338 0 42394 800
rect 42798 0 42854 800
rect 43258 0 43314 800
rect 43718 0 43774 800
rect 44178 0 44234 800
rect 44638 0 44694 800
rect 45098 0 45154 800
rect 45558 0 45614 800
rect 46018 0 46074 800
rect 46400 746 46428 1294
rect 46480 1284 46532 1290
rect 46480 1226 46532 1232
rect 46492 800 46520 1226
rect 47412 800 47440 2790
rect 47676 2372 47728 2378
rect 47676 2314 47728 2320
rect 47688 1766 47716 2314
rect 47860 1896 47912 1902
rect 47860 1838 47912 1844
rect 47676 1760 47728 1766
rect 47676 1702 47728 1708
rect 47872 800 47900 1838
rect 48332 1290 48360 3606
rect 48964 3528 49016 3534
rect 48964 3470 49016 3476
rect 48976 3194 49004 3470
rect 48964 3188 49016 3194
rect 48964 3130 49016 3136
rect 48872 3052 48924 3058
rect 48872 2994 48924 3000
rect 48780 2984 48832 2990
rect 48780 2926 48832 2932
rect 48792 2650 48820 2926
rect 48780 2644 48832 2650
rect 48780 2586 48832 2592
rect 48504 2304 48556 2310
rect 48504 2246 48556 2252
rect 48516 1426 48544 2246
rect 48504 1420 48556 1426
rect 48504 1362 48556 1368
rect 48884 1306 48912 2994
rect 49332 2984 49384 2990
rect 49332 2926 49384 2932
rect 49344 1358 49372 2926
rect 49528 2650 49556 3862
rect 49608 3732 49660 3738
rect 49608 3674 49660 3680
rect 49516 2644 49568 2650
rect 49516 2586 49568 2592
rect 49424 2440 49476 2446
rect 49424 2382 49476 2388
rect 49436 2038 49464 2382
rect 49424 2032 49476 2038
rect 49424 1974 49476 1980
rect 49620 1970 49648 3674
rect 49804 2514 49832 5102
rect 49884 3596 49936 3602
rect 49884 3538 49936 3544
rect 49792 2508 49844 2514
rect 49792 2450 49844 2456
rect 49896 1970 49924 3538
rect 49976 3392 50028 3398
rect 49976 3334 50028 3340
rect 49988 2514 50016 3334
rect 49976 2508 50028 2514
rect 49976 2450 50028 2456
rect 50172 2378 50200 5102
rect 50816 3942 50844 5646
rect 51264 5160 51316 5166
rect 51262 5128 51264 5137
rect 51356 5160 51408 5166
rect 51316 5128 51318 5137
rect 51356 5102 51408 5108
rect 51262 5063 51318 5072
rect 50804 3936 50856 3942
rect 50804 3878 50856 3884
rect 50712 3528 50764 3534
rect 50712 3470 50764 3476
rect 50436 3392 50488 3398
rect 50436 3334 50488 3340
rect 50448 3058 50476 3334
rect 50436 3052 50488 3058
rect 50436 2994 50488 3000
rect 50724 2650 50752 3470
rect 51368 3126 51396 5102
rect 51552 4010 51580 5646
rect 51724 5160 51776 5166
rect 51724 5102 51776 5108
rect 51736 4486 51764 5102
rect 51836 4922 52188 5972
rect 52460 5704 52512 5710
rect 52460 5646 52512 5652
rect 53840 5704 53892 5710
rect 53840 5646 53892 5652
rect 51836 4870 51858 4922
rect 51910 4870 51922 4922
rect 51974 4870 51986 4922
rect 52038 4870 52050 4922
rect 52102 4870 52114 4922
rect 52166 4870 52188 4922
rect 51724 4480 51776 4486
rect 51724 4422 51776 4428
rect 51540 4004 51592 4010
rect 51540 3946 51592 3952
rect 51836 3834 52188 4870
rect 52276 4004 52328 4010
rect 52276 3946 52328 3952
rect 51836 3782 51858 3834
rect 51910 3782 51922 3834
rect 51974 3782 51986 3834
rect 52038 3782 52050 3834
rect 52102 3782 52114 3834
rect 52166 3782 52188 3834
rect 51540 3460 51592 3466
rect 51540 3402 51592 3408
rect 51448 3392 51500 3398
rect 51448 3334 51500 3340
rect 51356 3120 51408 3126
rect 51356 3062 51408 3068
rect 51356 2916 51408 2922
rect 51356 2858 51408 2864
rect 51080 2848 51132 2854
rect 51080 2790 51132 2796
rect 51172 2848 51224 2854
rect 51172 2790 51224 2796
rect 50712 2644 50764 2650
rect 50712 2586 50764 2592
rect 51092 2514 51120 2790
rect 51080 2508 51132 2514
rect 51080 2450 51132 2456
rect 50160 2372 50212 2378
rect 50160 2314 50212 2320
rect 51184 2038 51212 2790
rect 51368 2446 51396 2858
rect 51460 2446 51488 3334
rect 51552 2650 51580 3402
rect 51724 3052 51776 3058
rect 51724 2994 51776 3000
rect 51632 2984 51684 2990
rect 51632 2926 51684 2932
rect 51540 2644 51592 2650
rect 51540 2586 51592 2592
rect 51356 2440 51408 2446
rect 51356 2382 51408 2388
rect 51448 2440 51500 2446
rect 51448 2382 51500 2388
rect 51172 2032 51224 2038
rect 51172 1974 51224 1980
rect 49608 1964 49660 1970
rect 49608 1906 49660 1912
rect 49884 1964 49936 1970
rect 49884 1906 49936 1912
rect 50620 1896 50672 1902
rect 50620 1838 50672 1844
rect 48320 1284 48372 1290
rect 48320 1226 48372 1232
rect 48792 1278 48912 1306
rect 49056 1352 49108 1358
rect 49056 1294 49108 1300
rect 49332 1352 49384 1358
rect 49332 1294 49384 1300
rect 48792 800 48820 1278
rect 49068 950 49096 1294
rect 49240 1284 49292 1290
rect 49240 1226 49292 1232
rect 49056 944 49108 950
rect 49056 886 49108 892
rect 49252 800 49280 1226
rect 50160 1216 50212 1222
rect 50160 1158 50212 1164
rect 50172 800 50200 1158
rect 50632 800 50660 1838
rect 51644 1358 51672 2926
rect 51448 1352 51500 1358
rect 51448 1294 51500 1300
rect 51632 1352 51684 1358
rect 51632 1294 51684 1300
rect 46388 740 46440 746
rect 46388 682 46440 688
rect 46478 0 46534 800
rect 46938 0 46994 800
rect 47398 0 47454 800
rect 47858 0 47914 800
rect 48318 0 48374 800
rect 48778 0 48834 800
rect 49238 0 49294 800
rect 49698 0 49754 800
rect 50158 0 50214 800
rect 50618 0 50674 800
rect 51078 0 51134 800
rect 51460 338 51488 1294
rect 51736 1170 51764 2994
rect 51552 1142 51764 1170
rect 51836 2746 52188 3782
rect 51836 2694 51858 2746
rect 51910 2694 51922 2746
rect 51974 2694 51986 2746
rect 52038 2694 52050 2746
rect 52102 2694 52114 2746
rect 52166 2694 52188 2746
rect 51836 2236 52188 2694
rect 51836 2180 51864 2236
rect 51920 2180 51944 2236
rect 52000 2180 52024 2236
rect 52080 2180 52104 2236
rect 52160 2180 52188 2236
rect 51836 2156 52188 2180
rect 51836 2100 51864 2156
rect 51920 2100 51944 2156
rect 52000 2100 52024 2156
rect 52080 2100 52104 2156
rect 52160 2100 52188 2156
rect 51836 2076 52188 2100
rect 51836 2020 51864 2076
rect 51920 2020 51944 2076
rect 52000 2020 52024 2076
rect 52080 2020 52104 2076
rect 52160 2020 52188 2076
rect 51836 1996 52188 2020
rect 51836 1940 51864 1996
rect 51920 1940 51944 1996
rect 52000 1940 52024 1996
rect 52080 1940 52104 1996
rect 52160 1940 52188 1996
rect 52288 1970 52316 3946
rect 52368 3392 52420 3398
rect 52368 3334 52420 3340
rect 52380 3126 52408 3334
rect 52368 3120 52420 3126
rect 52368 3062 52420 3068
rect 52472 2038 52500 5646
rect 53472 5364 53524 5370
rect 53472 5306 53524 5312
rect 52826 5264 52882 5273
rect 52826 5199 52828 5208
rect 52880 5199 52882 5208
rect 52828 5170 52880 5176
rect 53484 5166 53512 5306
rect 53288 5160 53340 5166
rect 53288 5102 53340 5108
rect 53380 5160 53432 5166
rect 53380 5102 53432 5108
rect 53472 5160 53524 5166
rect 53472 5102 53524 5108
rect 53300 4622 53328 5102
rect 53288 4616 53340 4622
rect 53288 4558 53340 4564
rect 53392 4162 53420 5102
rect 53300 4146 53420 4162
rect 53288 4140 53420 4146
rect 53340 4134 53420 4140
rect 53288 4082 53340 4088
rect 52644 3528 52696 3534
rect 52644 3470 52696 3476
rect 53012 3528 53064 3534
rect 53012 3470 53064 3476
rect 52656 3194 52684 3470
rect 52644 3188 52696 3194
rect 52644 3130 52696 3136
rect 52644 2984 52696 2990
rect 52644 2926 52696 2932
rect 52656 2038 52684 2926
rect 52920 2916 52972 2922
rect 52920 2858 52972 2864
rect 52460 2032 52512 2038
rect 52460 1974 52512 1980
rect 52644 2032 52696 2038
rect 52644 1974 52696 1980
rect 51836 1658 52188 1940
rect 52276 1964 52328 1970
rect 52276 1906 52328 1912
rect 51836 1606 51858 1658
rect 51910 1606 51922 1658
rect 51974 1606 51986 1658
rect 52038 1606 52050 1658
rect 52102 1606 52114 1658
rect 52166 1606 52188 1658
rect 51552 800 51580 1142
rect 51836 1040 52188 1606
rect 52368 1284 52420 1290
rect 52368 1226 52420 1232
rect 52012 870 52132 898
rect 52012 800 52040 870
rect 51448 332 51500 338
rect 51448 274 51500 280
rect 51538 0 51594 800
rect 51998 0 52054 800
rect 52104 762 52132 870
rect 52380 762 52408 1226
rect 52932 800 52960 2858
rect 53024 2650 53052 3470
rect 53852 3126 53880 5646
rect 54188 5466 54540 5944
rect 55048 5710 55076 7210
rect 58624 7064 58676 7070
rect 58624 7006 58676 7012
rect 56508 6860 56560 6866
rect 56508 6802 56560 6808
rect 55772 6792 55824 6798
rect 55824 6740 55996 6746
rect 55772 6734 55996 6740
rect 55784 6718 55996 6734
rect 55968 6662 55996 6718
rect 55956 6656 56008 6662
rect 55956 6598 56008 6604
rect 56324 6180 56376 6186
rect 56324 6122 56376 6128
rect 56232 6112 56284 6118
rect 56232 6054 56284 6060
rect 55036 5704 55088 5710
rect 55036 5646 55088 5652
rect 54188 5414 54210 5466
rect 54262 5414 54274 5466
rect 54326 5414 54338 5466
rect 54390 5414 54402 5466
rect 54454 5414 54466 5466
rect 54518 5414 54540 5466
rect 54024 5364 54076 5370
rect 54024 5306 54076 5312
rect 54036 4826 54064 5306
rect 54024 4820 54076 4826
rect 54024 4762 54076 4768
rect 54188 4588 54540 5414
rect 55864 5296 55916 5302
rect 55864 5238 55916 5244
rect 54852 5160 54904 5166
rect 54850 5128 54852 5137
rect 55404 5160 55456 5166
rect 54904 5128 54906 5137
rect 55404 5102 55456 5108
rect 54850 5063 54906 5072
rect 54188 4532 54216 4588
rect 54272 4532 54296 4588
rect 54352 4532 54376 4588
rect 54432 4532 54456 4588
rect 54512 4532 54540 4588
rect 54188 4508 54540 4532
rect 54188 4452 54216 4508
rect 54272 4452 54296 4508
rect 54352 4452 54376 4508
rect 54432 4452 54456 4508
rect 54512 4452 54540 4508
rect 54188 4428 54540 4452
rect 54188 4378 54216 4428
rect 54272 4378 54296 4428
rect 54352 4378 54376 4428
rect 54432 4378 54456 4428
rect 54512 4378 54540 4428
rect 54188 4326 54210 4378
rect 54272 4372 54274 4378
rect 54454 4372 54456 4378
rect 54262 4348 54274 4372
rect 54326 4348 54338 4372
rect 54390 4348 54402 4372
rect 54454 4348 54466 4372
rect 54272 4326 54274 4348
rect 54454 4326 54456 4348
rect 54518 4326 54540 4378
rect 54188 4292 54216 4326
rect 54272 4292 54296 4326
rect 54352 4292 54376 4326
rect 54432 4292 54456 4326
rect 54512 4292 54540 4326
rect 53932 3596 53984 3602
rect 53932 3538 53984 3544
rect 53840 3120 53892 3126
rect 53840 3062 53892 3068
rect 53012 2644 53064 2650
rect 53012 2586 53064 2592
rect 53196 2304 53248 2310
rect 53196 2246 53248 2252
rect 53208 1970 53236 2246
rect 53196 1964 53248 1970
rect 53196 1906 53248 1912
rect 53380 1896 53432 1902
rect 53380 1838 53432 1844
rect 53392 800 53420 1838
rect 53944 1222 53972 3538
rect 54024 3460 54076 3466
rect 54024 3402 54076 3408
rect 54036 2514 54064 3402
rect 54188 3290 54540 4292
rect 55416 4214 55444 5102
rect 55496 5024 55548 5030
rect 55496 4966 55548 4972
rect 55508 4214 55536 4966
rect 55404 4208 55456 4214
rect 55404 4150 55456 4156
rect 55496 4208 55548 4214
rect 55496 4150 55548 4156
rect 55876 4146 55904 5238
rect 56244 5030 56272 6054
rect 56336 5710 56364 6122
rect 56324 5704 56376 5710
rect 56324 5646 56376 5652
rect 56232 5024 56284 5030
rect 56232 4966 56284 4972
rect 56416 5024 56468 5030
rect 56416 4966 56468 4972
rect 56428 4282 56456 4966
rect 56416 4276 56468 4282
rect 56416 4218 56468 4224
rect 55864 4140 55916 4146
rect 55864 4082 55916 4088
rect 55864 3936 55916 3942
rect 55864 3878 55916 3884
rect 55876 3738 55904 3878
rect 55864 3732 55916 3738
rect 55864 3674 55916 3680
rect 54668 3664 54720 3670
rect 54668 3606 54720 3612
rect 54188 3238 54210 3290
rect 54262 3238 54274 3290
rect 54326 3238 54338 3290
rect 54390 3238 54402 3290
rect 54454 3238 54466 3290
rect 54518 3238 54540 3290
rect 54024 2508 54076 2514
rect 54024 2450 54076 2456
rect 54188 2202 54540 3238
rect 54576 2984 54628 2990
rect 54576 2926 54628 2932
rect 54188 2150 54210 2202
rect 54262 2150 54274 2202
rect 54326 2150 54338 2202
rect 54390 2150 54402 2202
rect 54454 2150 54466 2202
rect 54518 2150 54540 2202
rect 54024 1352 54076 1358
rect 54024 1294 54076 1300
rect 53932 1216 53984 1222
rect 53932 1158 53984 1164
rect 52104 734 52408 762
rect 52458 0 52514 800
rect 52918 0 52974 800
rect 53378 0 53434 800
rect 53838 0 53894 800
rect 54036 542 54064 1294
rect 54188 1114 54540 2150
rect 54188 1062 54210 1114
rect 54262 1062 54274 1114
rect 54326 1062 54338 1114
rect 54390 1062 54402 1114
rect 54454 1062 54466 1114
rect 54518 1062 54540 1114
rect 54188 1040 54540 1062
rect 54312 870 54432 898
rect 54312 800 54340 870
rect 54024 536 54076 542
rect 54024 478 54076 484
rect 54298 0 54354 800
rect 54404 762 54432 870
rect 54588 762 54616 2926
rect 54680 2582 54708 3606
rect 55956 3528 56008 3534
rect 55956 3470 56008 3476
rect 55588 3392 55640 3398
rect 55588 3334 55640 3340
rect 55600 3058 55628 3334
rect 54944 3052 54996 3058
rect 54944 2994 54996 3000
rect 55588 3052 55640 3058
rect 55588 2994 55640 3000
rect 54668 2576 54720 2582
rect 54668 2518 54720 2524
rect 54956 1970 54984 2994
rect 55680 2984 55732 2990
rect 55680 2926 55732 2932
rect 55312 2916 55364 2922
rect 55312 2858 55364 2864
rect 55220 2848 55272 2854
rect 55220 2790 55272 2796
rect 55232 2514 55260 2790
rect 55220 2508 55272 2514
rect 55220 2450 55272 2456
rect 55324 1970 55352 2858
rect 54944 1964 54996 1970
rect 54944 1906 54996 1912
rect 55312 1964 55364 1970
rect 55312 1906 55364 1912
rect 54760 1284 54812 1290
rect 54760 1226 54812 1232
rect 54772 800 54800 1226
rect 55692 800 55720 2926
rect 55968 2582 55996 3470
rect 55956 2576 56008 2582
rect 55956 2518 56008 2524
rect 56048 2304 56100 2310
rect 56048 2246 56100 2252
rect 55864 2100 55916 2106
rect 55864 2042 55916 2048
rect 55876 1426 55904 2042
rect 56060 1970 56088 2246
rect 56520 2106 56548 6802
rect 58530 6352 58586 6361
rect 58530 6287 58586 6296
rect 57610 6216 57666 6225
rect 57610 6151 57666 6160
rect 56692 5704 56744 5710
rect 56692 5646 56744 5652
rect 56598 5264 56654 5273
rect 56598 5199 56600 5208
rect 56652 5199 56654 5208
rect 56600 5170 56652 5176
rect 56704 4486 56732 5646
rect 56692 4480 56744 4486
rect 56692 4422 56744 4428
rect 57060 2984 57112 2990
rect 57060 2926 57112 2932
rect 56600 2916 56652 2922
rect 56600 2858 56652 2864
rect 56612 2514 56640 2858
rect 56876 2848 56928 2854
rect 56876 2790 56928 2796
rect 56968 2848 57020 2854
rect 56968 2790 57020 2796
rect 56888 2514 56916 2790
rect 56600 2508 56652 2514
rect 56600 2450 56652 2456
rect 56876 2508 56928 2514
rect 56876 2450 56928 2456
rect 56692 2440 56744 2446
rect 56692 2382 56744 2388
rect 56508 2100 56560 2106
rect 56508 2042 56560 2048
rect 56048 1964 56100 1970
rect 56048 1906 56100 1912
rect 56140 1896 56192 1902
rect 56140 1838 56192 1844
rect 55864 1420 55916 1426
rect 55864 1362 55916 1368
rect 56152 800 56180 1838
rect 56704 1358 56732 2382
rect 56980 1902 57008 2790
rect 56968 1896 57020 1902
rect 56968 1838 57020 1844
rect 56692 1352 56744 1358
rect 56692 1294 56744 1300
rect 57072 800 57100 2926
rect 57244 2372 57296 2378
rect 57244 2314 57296 2320
rect 57256 1358 57284 2314
rect 57624 1970 57652 6151
rect 58544 5574 58572 6287
rect 58532 5568 58584 5574
rect 58532 5510 58584 5516
rect 58636 4010 58664 7006
rect 61476 6928 61528 6934
rect 61476 6870 61528 6876
rect 60924 6656 60976 6662
rect 60922 6624 60924 6633
rect 61108 6656 61160 6662
rect 60976 6624 60978 6633
rect 61108 6598 61160 6604
rect 61382 6624 61438 6633
rect 60922 6559 60978 6568
rect 61120 6390 61148 6598
rect 61382 6559 61438 6568
rect 61108 6384 61160 6390
rect 61108 6326 61160 6332
rect 61108 5908 61160 5914
rect 61108 5850 61160 5856
rect 61120 5794 61148 5850
rect 60280 5772 60332 5778
rect 60464 5772 60516 5778
rect 60280 5714 60332 5720
rect 60384 5732 60464 5760
rect 60292 5642 60320 5714
rect 60280 5636 60332 5642
rect 60280 5578 60332 5584
rect 60384 5370 60412 5732
rect 60464 5714 60516 5720
rect 60660 5766 61148 5794
rect 61396 5778 61424 6559
rect 61292 5772 61344 5778
rect 60372 5364 60424 5370
rect 60372 5306 60424 5312
rect 60556 5296 60608 5302
rect 60556 5238 60608 5244
rect 60568 4622 60596 5238
rect 60556 4616 60608 4622
rect 60556 4558 60608 4564
rect 60464 4276 60516 4282
rect 60464 4218 60516 4224
rect 58624 4004 58676 4010
rect 58624 3946 58676 3952
rect 59084 3664 59136 3670
rect 59084 3606 59136 3612
rect 58164 3392 58216 3398
rect 58164 3334 58216 3340
rect 58176 3058 58204 3334
rect 58164 3052 58216 3058
rect 58164 2994 58216 3000
rect 58532 2916 58584 2922
rect 58532 2858 58584 2864
rect 58440 2440 58492 2446
rect 58440 2382 58492 2388
rect 58452 2106 58480 2382
rect 58440 2100 58492 2106
rect 58440 2042 58492 2048
rect 57612 1964 57664 1970
rect 57612 1906 57664 1912
rect 58544 1544 58572 2858
rect 58900 2848 58952 2854
rect 58900 2790 58952 2796
rect 58912 2514 58940 2790
rect 58900 2508 58952 2514
rect 58900 2450 58952 2456
rect 58900 1896 58952 1902
rect 58900 1838 58952 1844
rect 58452 1516 58572 1544
rect 57244 1352 57296 1358
rect 57244 1294 57296 1300
rect 57520 1284 57572 1290
rect 57520 1226 57572 1232
rect 57532 800 57560 1226
rect 58452 800 58480 1516
rect 58912 800 58940 1838
rect 59096 1358 59124 3606
rect 60372 3528 60424 3534
rect 60372 3470 60424 3476
rect 59176 3460 59228 3466
rect 59176 3402 59228 3408
rect 59188 3058 59216 3402
rect 59268 3120 59320 3126
rect 59268 3062 59320 3068
rect 59176 3052 59228 3058
rect 59176 2994 59228 3000
rect 59280 1358 59308 3062
rect 59820 2984 59872 2990
rect 59820 2926 59872 2932
rect 59728 2440 59780 2446
rect 59728 2382 59780 2388
rect 59452 2304 59504 2310
rect 59452 2246 59504 2252
rect 59544 2304 59596 2310
rect 59544 2246 59596 2252
rect 59464 1358 59492 2246
rect 59556 1902 59584 2246
rect 59544 1896 59596 1902
rect 59544 1838 59596 1844
rect 59740 1562 59768 2382
rect 59728 1556 59780 1562
rect 59728 1498 59780 1504
rect 59084 1352 59136 1358
rect 59084 1294 59136 1300
rect 59268 1352 59320 1358
rect 59268 1294 59320 1300
rect 59452 1352 59504 1358
rect 59452 1294 59504 1300
rect 59832 800 59860 2926
rect 59912 2848 59964 2854
rect 59912 2790 59964 2796
rect 59924 2514 59952 2790
rect 59912 2508 59964 2514
rect 59912 2450 59964 2456
rect 60384 2106 60412 3470
rect 60372 2100 60424 2106
rect 60372 2042 60424 2048
rect 60476 1970 60504 4218
rect 60660 2582 60688 5766
rect 61292 5714 61344 5720
rect 61384 5772 61436 5778
rect 61384 5714 61436 5720
rect 61304 5658 61332 5714
rect 61488 5658 61516 6870
rect 61304 5630 61516 5658
rect 61836 4922 62188 5972
rect 61836 4870 61858 4922
rect 61910 4870 61922 4922
rect 61974 4870 61986 4922
rect 62038 4870 62050 4922
rect 62102 4870 62114 4922
rect 62166 4870 62188 4922
rect 61836 3834 62188 4870
rect 61836 3782 61858 3834
rect 61910 3782 61922 3834
rect 61974 3782 61986 3834
rect 62038 3782 62050 3834
rect 62102 3782 62114 3834
rect 62166 3782 62188 3834
rect 60740 3460 60792 3466
rect 60740 3402 60792 3408
rect 60752 3194 60780 3402
rect 60740 3188 60792 3194
rect 60740 3130 60792 3136
rect 61384 2984 61436 2990
rect 61384 2926 61436 2932
rect 61568 2984 61620 2990
rect 61568 2926 61620 2932
rect 61108 2848 61160 2854
rect 61108 2790 61160 2796
rect 60648 2576 60700 2582
rect 60648 2518 60700 2524
rect 61120 2514 61148 2790
rect 61108 2508 61160 2514
rect 61108 2450 61160 2456
rect 61200 2304 61252 2310
rect 61200 2246 61252 2252
rect 61212 1970 61240 2246
rect 61396 2106 61424 2926
rect 61580 2582 61608 2926
rect 61836 2746 62188 3782
rect 61836 2694 61858 2746
rect 61910 2694 61922 2746
rect 61974 2694 61986 2746
rect 62038 2694 62050 2746
rect 62102 2694 62114 2746
rect 62166 2694 62188 2746
rect 61568 2576 61620 2582
rect 61568 2518 61620 2524
rect 61568 2440 61620 2446
rect 61568 2382 61620 2388
rect 61384 2100 61436 2106
rect 61384 2042 61436 2048
rect 60464 1964 60516 1970
rect 60464 1906 60516 1912
rect 61200 1964 61252 1970
rect 61200 1906 61252 1912
rect 60280 1284 60332 1290
rect 60280 1226 60332 1232
rect 60292 800 60320 1226
rect 61212 870 61332 898
rect 61212 800 61240 870
rect 54404 734 54616 762
rect 54758 0 54814 800
rect 55218 0 55274 800
rect 55678 0 55734 800
rect 56138 0 56194 800
rect 56598 0 56654 800
rect 57058 0 57114 800
rect 57518 0 57574 800
rect 57978 0 58034 800
rect 58438 0 58494 800
rect 58898 0 58954 800
rect 59358 0 59414 800
rect 59818 0 59874 800
rect 60278 0 60334 800
rect 60738 0 60794 800
rect 61198 0 61254 800
rect 61304 762 61332 870
rect 61580 762 61608 2382
rect 61660 2372 61712 2378
rect 61660 2314 61712 2320
rect 61672 1494 61700 2314
rect 61836 2236 62188 2694
rect 61836 2180 61864 2236
rect 61920 2180 61944 2236
rect 62000 2180 62024 2236
rect 62080 2180 62104 2236
rect 62160 2180 62188 2236
rect 61836 2156 62188 2180
rect 61836 2100 61864 2156
rect 61920 2100 61944 2156
rect 62000 2100 62024 2156
rect 62080 2100 62104 2156
rect 62160 2100 62188 2156
rect 61836 2076 62188 2100
rect 61836 2020 61864 2076
rect 61920 2020 61944 2076
rect 62000 2020 62024 2076
rect 62080 2020 62104 2076
rect 62160 2020 62188 2076
rect 61836 1996 62188 2020
rect 61836 1940 61864 1996
rect 61920 1940 61944 1996
rect 62000 1940 62024 1996
rect 62080 1940 62104 1996
rect 62160 1940 62188 1996
rect 61836 1658 62188 1940
rect 61836 1606 61858 1658
rect 61910 1606 61922 1658
rect 61974 1606 61986 1658
rect 62038 1606 62050 1658
rect 62102 1606 62114 1658
rect 62166 1606 62188 1658
rect 61660 1488 61712 1494
rect 61660 1430 61712 1436
rect 61660 1284 61712 1290
rect 61660 1226 61712 1232
rect 61672 800 61700 1226
rect 61836 1040 62188 1606
rect 62316 1358 62344 7278
rect 62684 5953 62712 7346
rect 62764 7200 62816 7206
rect 62764 7142 62816 7148
rect 62776 6594 62804 7142
rect 62764 6588 62816 6594
rect 62764 6530 62816 6536
rect 63144 6526 63172 7414
rect 63132 6520 63184 6526
rect 63132 6462 63184 6468
rect 62670 5944 62726 5953
rect 62670 5879 62726 5888
rect 63236 5030 63264 7822
rect 63420 7818 63448 11086
rect 63500 10344 63552 10350
rect 63500 10286 63552 10292
rect 63408 7812 63460 7818
rect 63408 7754 63460 7760
rect 63316 6996 63368 7002
rect 63316 6938 63368 6944
rect 63328 6254 63356 6938
rect 63512 6934 63540 10286
rect 63604 7614 63632 11206
rect 63592 7608 63644 7614
rect 63592 7550 63644 7556
rect 63500 6928 63552 6934
rect 63500 6870 63552 6876
rect 63316 6248 63368 6254
rect 63316 6190 63368 6196
rect 63592 6248 63644 6254
rect 63592 6190 63644 6196
rect 63224 5024 63276 5030
rect 63224 4966 63276 4972
rect 63604 3670 63632 6190
rect 63592 3664 63644 3670
rect 63592 3606 63644 3612
rect 63408 3052 63460 3058
rect 63408 2994 63460 3000
rect 63316 2984 63368 2990
rect 63316 2926 63368 2932
rect 62580 2916 62632 2922
rect 62580 2858 62632 2864
rect 62592 2514 62620 2858
rect 63328 2582 63356 2926
rect 63316 2576 63368 2582
rect 63316 2518 63368 2524
rect 62580 2508 62632 2514
rect 62580 2450 62632 2456
rect 62672 2508 62724 2514
rect 62672 2450 62724 2456
rect 62488 2304 62540 2310
rect 62488 2246 62540 2252
rect 62500 1970 62528 2246
rect 62488 1964 62540 1970
rect 62488 1906 62540 1912
rect 62684 1902 62712 2450
rect 62764 2440 62816 2446
rect 62764 2382 62816 2388
rect 62672 1896 62724 1902
rect 62672 1838 62724 1844
rect 62396 1828 62448 1834
rect 62396 1770 62448 1776
rect 62408 1358 62436 1770
rect 62304 1352 62356 1358
rect 62304 1294 62356 1300
rect 62396 1352 62448 1358
rect 62396 1294 62448 1300
rect 62776 1272 62804 2382
rect 63040 1896 63092 1902
rect 63040 1838 63092 1844
rect 62592 1244 62804 1272
rect 62592 800 62620 1244
rect 63052 800 63080 1838
rect 63420 1358 63448 2994
rect 63132 1352 63184 1358
rect 63132 1294 63184 1300
rect 63408 1352 63460 1358
rect 63408 1294 63460 1300
rect 61304 734 61608 762
rect 61658 0 61714 800
rect 62118 0 62174 800
rect 62578 0 62634 800
rect 63038 0 63094 800
rect 63144 406 63172 1294
rect 63696 1222 63724 56578
rect 63776 52488 63828 52494
rect 63776 52430 63828 52436
rect 63684 1216 63736 1222
rect 63684 1158 63736 1164
rect 63132 400 63184 406
rect 63132 342 63184 348
rect 63498 0 63554 800
rect 63788 542 63816 52430
rect 63868 50312 63920 50318
rect 63868 50254 63920 50260
rect 63880 11490 63908 50254
rect 63960 43172 64012 43178
rect 63960 43114 64012 43120
rect 63868 11484 63920 11490
rect 63868 11426 63920 11432
rect 63868 11348 63920 11354
rect 63868 11290 63920 11296
rect 63880 4282 63908 11290
rect 63868 4276 63920 4282
rect 63868 4218 63920 4224
rect 63972 1952 64000 43114
rect 64052 40996 64104 41002
rect 64052 40938 64104 40944
rect 63880 1924 64000 1952
rect 63880 1766 63908 1924
rect 63960 1828 64012 1834
rect 63960 1770 64012 1776
rect 63868 1760 63920 1766
rect 63868 1702 63920 1708
rect 63972 800 64000 1770
rect 64064 814 64092 40938
rect 64144 35692 64196 35698
rect 64144 35634 64196 35640
rect 64156 6089 64184 35634
rect 64236 27532 64288 27538
rect 64236 27474 64288 27480
rect 64248 7274 64276 27474
rect 64328 26988 64380 26994
rect 64328 26930 64380 26936
rect 64340 16574 64368 26930
rect 64340 16546 64460 16574
rect 64328 11416 64380 11422
rect 64328 11358 64380 11364
rect 64236 7268 64288 7274
rect 64236 7210 64288 7216
rect 64340 6254 64368 11358
rect 64328 6248 64380 6254
rect 64328 6190 64380 6196
rect 64432 6089 64460 16546
rect 64512 11484 64564 11490
rect 64512 11426 64564 11432
rect 64524 7070 64552 11426
rect 64512 7064 64564 7070
rect 64512 7006 64564 7012
rect 64142 6080 64198 6089
rect 64142 6015 64198 6024
rect 64418 6080 64474 6089
rect 64418 6015 64474 6024
rect 64188 5466 64540 5972
rect 64188 5414 64210 5466
rect 64262 5414 64274 5466
rect 64326 5414 64338 5466
rect 64390 5414 64402 5466
rect 64454 5414 64466 5466
rect 64518 5414 64540 5466
rect 64188 4588 64540 5414
rect 64188 4532 64216 4588
rect 64272 4532 64296 4588
rect 64352 4532 64376 4588
rect 64432 4532 64456 4588
rect 64512 4532 64540 4588
rect 64188 4508 64540 4532
rect 64188 4452 64216 4508
rect 64272 4452 64296 4508
rect 64352 4452 64376 4508
rect 64432 4452 64456 4508
rect 64512 4452 64540 4508
rect 64188 4428 64540 4452
rect 64188 4378 64216 4428
rect 64272 4378 64296 4428
rect 64352 4378 64376 4428
rect 64432 4378 64456 4428
rect 64512 4378 64540 4428
rect 64188 4326 64210 4378
rect 64272 4372 64274 4378
rect 64454 4372 64456 4378
rect 64262 4348 64274 4372
rect 64326 4348 64338 4372
rect 64390 4348 64402 4372
rect 64454 4348 64466 4372
rect 64272 4326 64274 4348
rect 64454 4326 64456 4348
rect 64518 4326 64540 4378
rect 64188 4292 64216 4326
rect 64272 4292 64296 4326
rect 64352 4292 64376 4326
rect 64432 4292 64456 4326
rect 64512 4292 64540 4326
rect 64188 3290 64540 4292
rect 64188 3238 64210 3290
rect 64262 3238 64274 3290
rect 64326 3238 64338 3290
rect 64390 3238 64402 3290
rect 64454 3238 64466 3290
rect 64518 3238 64540 3290
rect 64188 2202 64540 3238
rect 64188 2150 64210 2202
rect 64262 2150 64274 2202
rect 64326 2150 64338 2202
rect 64390 2150 64402 2202
rect 64454 2150 64466 2202
rect 64518 2150 64540 2202
rect 64188 1114 64540 2150
rect 64616 1970 64644 71742
rect 64892 71126 64920 73170
rect 65156 72208 65208 72214
rect 65156 72150 65208 72156
rect 64880 71120 64932 71126
rect 64880 71062 64932 71068
rect 64892 68950 64920 71062
rect 64880 68944 64932 68950
rect 64880 68886 64932 68892
rect 65064 67856 65116 67862
rect 65064 67798 65116 67804
rect 64880 66496 64932 66502
rect 64880 66438 64932 66444
rect 64892 64326 64920 66438
rect 64880 64320 64932 64326
rect 64880 64262 64932 64268
rect 64892 62150 64920 64262
rect 64972 63572 65024 63578
rect 64972 63514 65024 63520
rect 64880 62144 64932 62150
rect 64880 62086 64932 62092
rect 64892 60246 64920 62086
rect 64880 60240 64932 60246
rect 64880 60182 64932 60188
rect 64892 58070 64920 60182
rect 64880 58064 64932 58070
rect 64880 58006 64932 58012
rect 64892 55622 64920 58006
rect 64880 55616 64932 55622
rect 64880 55558 64932 55564
rect 64892 53582 64920 55558
rect 64880 53576 64932 53582
rect 64880 53518 64932 53524
rect 64892 51542 64920 53518
rect 64880 51536 64932 51542
rect 64880 51478 64932 51484
rect 64984 48890 65012 63514
rect 65076 52018 65104 67798
rect 65168 55418 65196 72150
rect 65248 70032 65300 70038
rect 65248 69974 65300 69980
rect 65156 55412 65208 55418
rect 65156 55354 65208 55360
rect 65260 53242 65288 69974
rect 65352 58682 65380 76502
rect 65432 74656 65484 74662
rect 65432 74598 65484 74604
rect 65340 58676 65392 58682
rect 65340 58618 65392 58624
rect 65444 57050 65472 74598
rect 65536 61946 65564 80922
rect 65616 78736 65668 78742
rect 65616 78678 65668 78684
rect 65524 61940 65576 61946
rect 65524 61882 65576 61888
rect 65628 60314 65656 78678
rect 65720 63510 65748 83098
rect 71688 83020 71740 83026
rect 71688 82962 71740 82968
rect 70676 80844 70728 80850
rect 70676 80786 70728 80792
rect 68652 78668 68704 78674
rect 68652 78610 68704 78616
rect 68100 76492 68152 76498
rect 68100 76434 68152 76440
rect 65892 74112 65944 74118
rect 65892 74054 65944 74060
rect 65800 68944 65852 68950
rect 65800 68886 65852 68892
rect 65708 63504 65760 63510
rect 65708 63446 65760 63452
rect 65616 60308 65668 60314
rect 65616 60250 65668 60256
rect 65708 59152 65760 59158
rect 65708 59094 65760 59100
rect 65432 57044 65484 57050
rect 65432 56986 65484 56992
rect 65524 56976 65576 56982
rect 65524 56918 65576 56924
rect 65340 54800 65392 54806
rect 65340 54742 65392 54748
rect 65248 53236 65300 53242
rect 65248 53178 65300 53184
rect 65064 52012 65116 52018
rect 65064 51954 65116 51960
rect 65156 50448 65208 50454
rect 65156 50390 65208 50396
rect 64972 48884 65024 48890
rect 64972 48826 65024 48832
rect 64972 47728 65024 47734
rect 64972 47670 65024 47676
rect 64880 47388 64932 47394
rect 64880 47330 64932 47336
rect 64892 36378 64920 47330
rect 64984 44742 65012 47670
rect 65064 45960 65116 45966
rect 65064 45902 65116 45908
rect 64972 44736 65024 44742
rect 64972 44678 65024 44684
rect 64972 44600 65024 44606
rect 64972 44542 65024 44548
rect 64984 36786 65012 44542
rect 64972 36780 65024 36786
rect 64972 36722 65024 36728
rect 64972 36576 65024 36582
rect 64972 36518 65024 36524
rect 64880 36372 64932 36378
rect 64880 36314 64932 36320
rect 64880 35216 64932 35222
rect 64880 35158 64932 35164
rect 64892 33318 64920 35158
rect 64880 33312 64932 33318
rect 64880 33254 64932 33260
rect 64892 31142 64920 33254
rect 64880 31136 64932 31142
rect 64880 31078 64932 31084
rect 64892 28694 64920 31078
rect 64880 28688 64932 28694
rect 64880 28630 64932 28636
rect 64892 26790 64920 28630
rect 64880 26784 64932 26790
rect 64880 26726 64932 26732
rect 64880 24336 64932 24342
rect 64880 24278 64932 24284
rect 64892 23730 64920 24278
rect 64880 23724 64932 23730
rect 64880 23666 64932 23672
rect 64880 23520 64932 23526
rect 64880 23462 64932 23468
rect 64788 21344 64840 21350
rect 64788 21286 64840 21292
rect 64696 16108 64748 16114
rect 64696 16050 64748 16056
rect 64708 3670 64736 16050
rect 64696 3664 64748 3670
rect 64696 3606 64748 3612
rect 64696 3528 64748 3534
rect 64696 3470 64748 3476
rect 64708 2582 64736 3470
rect 64696 2576 64748 2582
rect 64696 2518 64748 2524
rect 64800 2378 64828 21286
rect 64892 18290 64920 23462
rect 64880 18284 64932 18290
rect 64880 18226 64932 18232
rect 64880 16652 64932 16658
rect 64880 16594 64932 16600
rect 64892 13530 64920 16594
rect 64880 13524 64932 13530
rect 64880 13466 64932 13472
rect 64880 13388 64932 13394
rect 64880 13330 64932 13336
rect 64892 11370 64920 13330
rect 64984 11558 65012 36518
rect 65076 34746 65104 45902
rect 65168 42106 65196 50390
rect 65352 42362 65380 54742
rect 65432 52624 65484 52630
rect 65432 52566 65484 52572
rect 65340 42356 65392 42362
rect 65340 42298 65392 42304
rect 65168 42078 65288 42106
rect 65444 42090 65472 52566
rect 65536 43994 65564 56918
rect 65616 52488 65668 52494
rect 65616 52430 65668 52436
rect 65628 52154 65656 52430
rect 65616 52148 65668 52154
rect 65616 52090 65668 52096
rect 65720 51074 65748 59094
rect 65812 53650 65840 68886
rect 65800 53644 65852 53650
rect 65800 53586 65852 53592
rect 65800 51536 65852 51542
rect 65800 51478 65852 51484
rect 65628 51046 65748 51074
rect 65628 45558 65656 51046
rect 65812 46186 65840 51478
rect 65720 46158 65840 46186
rect 65616 45552 65668 45558
rect 65616 45494 65668 45500
rect 65616 44736 65668 44742
rect 65616 44678 65668 44684
rect 65524 43988 65576 43994
rect 65524 43930 65576 43936
rect 65156 41744 65208 41750
rect 65156 41686 65208 41692
rect 65168 39846 65196 41686
rect 65156 39840 65208 39846
rect 65156 39782 65208 39788
rect 65168 37398 65196 39782
rect 65260 39098 65288 42078
rect 65432 42084 65484 42090
rect 65432 42026 65484 42032
rect 65432 41812 65484 41818
rect 65432 41754 65484 41760
rect 65340 40588 65392 40594
rect 65340 40530 65392 40536
rect 65248 39092 65300 39098
rect 65248 39034 65300 39040
rect 65156 37392 65208 37398
rect 65156 37334 65208 37340
rect 65168 35222 65196 37334
rect 65156 35216 65208 35222
rect 65156 35158 65208 35164
rect 65064 34740 65116 34746
rect 65064 34682 65116 34688
rect 65064 34536 65116 34542
rect 65064 34478 65116 34484
rect 64972 11552 65024 11558
rect 64972 11494 65024 11500
rect 64892 11342 65012 11370
rect 64984 11286 65012 11342
rect 64972 11280 65024 11286
rect 64972 11222 65024 11228
rect 64880 10600 64932 10606
rect 64880 10542 64932 10548
rect 64892 7993 64920 10542
rect 64984 9382 65012 11222
rect 64972 9376 65024 9382
rect 64972 9318 65024 9324
rect 64878 7984 64934 7993
rect 64878 7919 64934 7928
rect 64880 7880 64932 7886
rect 64880 7822 64932 7828
rect 64788 2372 64840 2378
rect 64788 2314 64840 2320
rect 64604 1964 64656 1970
rect 64604 1906 64656 1912
rect 64788 1896 64840 1902
rect 64788 1838 64840 1844
rect 64188 1062 64210 1114
rect 64262 1062 64274 1114
rect 64326 1062 64338 1114
rect 64390 1062 64402 1114
rect 64454 1062 64466 1114
rect 64518 1062 64540 1114
rect 64188 1040 64540 1062
rect 64432 870 64552 898
rect 64052 808 64104 814
rect 63776 536 63828 542
rect 63776 478 63828 484
rect 63958 0 64014 800
rect 64432 800 64460 870
rect 64052 750 64104 756
rect 64418 0 64474 800
rect 64524 762 64552 870
rect 64800 762 64828 1838
rect 64892 898 64920 7822
rect 64984 6186 65012 9318
rect 64972 6180 65024 6186
rect 64972 6122 65024 6128
rect 64972 3528 65024 3534
rect 64972 3470 65024 3476
rect 64984 3126 65012 3470
rect 64972 3120 65024 3126
rect 64972 3062 65024 3068
rect 64972 2848 65024 2854
rect 64972 2790 65024 2796
rect 64984 2514 65012 2790
rect 64972 2508 65024 2514
rect 64972 2450 65024 2456
rect 64972 2304 65024 2310
rect 64972 2246 65024 2252
rect 64984 1426 65012 2246
rect 65076 1562 65104 34478
rect 65156 33992 65208 33998
rect 65156 33934 65208 33940
rect 65168 29034 65196 33934
rect 65248 32224 65300 32230
rect 65248 32166 65300 32172
rect 65156 29028 65208 29034
rect 65156 28970 65208 28976
rect 65156 27668 65208 27674
rect 65156 27610 65208 27616
rect 65168 21690 65196 27610
rect 65156 21684 65208 21690
rect 65156 21626 65208 21632
rect 65156 21412 65208 21418
rect 65156 21354 65208 21360
rect 65168 7886 65196 21354
rect 65156 7880 65208 7886
rect 65156 7822 65208 7828
rect 65156 7744 65208 7750
rect 65156 7686 65208 7692
rect 65064 1556 65116 1562
rect 65064 1498 65116 1504
rect 65168 1494 65196 7686
rect 65260 7562 65288 32166
rect 65352 31482 65380 40530
rect 65444 40186 65472 41754
rect 65432 40180 65484 40186
rect 65432 40122 65484 40128
rect 65524 39636 65576 39642
rect 65524 39578 65576 39584
rect 65432 38752 65484 38758
rect 65432 38694 65484 38700
rect 65340 31476 65392 31482
rect 65340 31418 65392 31424
rect 65444 30326 65472 38694
rect 65536 36922 65564 39578
rect 65628 37262 65656 44678
rect 65720 40594 65748 46158
rect 65800 44192 65852 44198
rect 65800 44134 65852 44140
rect 65812 41041 65840 44134
rect 65798 41032 65854 41041
rect 65798 40967 65854 40976
rect 65800 40928 65852 40934
rect 65800 40870 65852 40876
rect 65708 40588 65760 40594
rect 65708 40530 65760 40536
rect 65708 40384 65760 40390
rect 65708 40326 65760 40332
rect 65616 37256 65668 37262
rect 65616 37198 65668 37204
rect 65524 36916 65576 36922
rect 65524 36858 65576 36864
rect 65524 36780 65576 36786
rect 65524 36722 65576 36728
rect 65536 33658 65564 36722
rect 65616 35012 65668 35018
rect 65616 34954 65668 34960
rect 65524 33652 65576 33658
rect 65524 33594 65576 33600
rect 65432 30320 65484 30326
rect 65432 30262 65484 30268
rect 65340 30048 65392 30054
rect 65340 29990 65392 29996
rect 65352 7750 65380 29990
rect 65628 28762 65656 34954
rect 65720 34202 65748 40326
rect 65708 34196 65760 34202
rect 65708 34138 65760 34144
rect 65708 33448 65760 33454
rect 65708 33390 65760 33396
rect 65616 28756 65668 28762
rect 65616 28698 65668 28704
rect 65524 27872 65576 27878
rect 65524 27814 65576 27820
rect 65432 25696 65484 25702
rect 65432 25638 65484 25644
rect 65444 23225 65472 25638
rect 65430 23216 65486 23225
rect 65430 23151 65486 23160
rect 65432 23044 65484 23050
rect 65432 22986 65484 22992
rect 65444 18426 65472 22986
rect 65536 21418 65564 27814
rect 65616 24880 65668 24886
rect 65616 24822 65668 24828
rect 65628 23866 65656 24822
rect 65616 23860 65668 23866
rect 65616 23802 65668 23808
rect 65616 23724 65668 23730
rect 65616 23666 65668 23672
rect 65628 22658 65656 23666
rect 65720 22778 65748 33390
rect 65812 27470 65840 40870
rect 65800 27464 65852 27470
rect 65800 27406 65852 27412
rect 65708 22772 65760 22778
rect 65708 22714 65760 22720
rect 65628 22630 65748 22658
rect 65614 22536 65670 22545
rect 65614 22471 65670 22480
rect 65524 21412 65576 21418
rect 65524 21354 65576 21360
rect 65628 21298 65656 22471
rect 65720 22166 65748 22630
rect 65708 22160 65760 22166
rect 65708 22102 65760 22108
rect 65536 21270 65656 21298
rect 65536 19922 65564 21270
rect 65616 20936 65668 20942
rect 65616 20878 65668 20884
rect 65524 19916 65576 19922
rect 65524 19858 65576 19864
rect 65524 18760 65576 18766
rect 65524 18702 65576 18708
rect 65432 18420 65484 18426
rect 65432 18362 65484 18368
rect 65432 18284 65484 18290
rect 65432 18226 65484 18232
rect 65340 7744 65392 7750
rect 65340 7686 65392 7692
rect 65260 7534 65380 7562
rect 65246 7440 65302 7449
rect 65246 7375 65302 7384
rect 65260 3942 65288 7375
rect 65248 3936 65300 3942
rect 65248 3878 65300 3884
rect 65248 2984 65300 2990
rect 65248 2926 65300 2932
rect 65260 2650 65288 2926
rect 65248 2644 65300 2650
rect 65248 2586 65300 2592
rect 65352 2530 65380 7534
rect 65260 2502 65380 2530
rect 65156 1488 65208 1494
rect 65156 1430 65208 1436
rect 64972 1420 65024 1426
rect 64972 1362 65024 1368
rect 64892 870 65012 898
rect 64524 734 64828 762
rect 64878 0 64934 800
rect 64984 610 65012 870
rect 65260 678 65288 2502
rect 65340 2440 65392 2446
rect 65340 2382 65392 2388
rect 65352 800 65380 2382
rect 65444 882 65472 18226
rect 65536 14618 65564 18702
rect 65628 17338 65656 20878
rect 65720 20330 65748 22102
rect 65708 20324 65760 20330
rect 65708 20266 65760 20272
rect 65720 18086 65748 20266
rect 65708 18080 65760 18086
rect 65708 18022 65760 18028
rect 65616 17332 65668 17338
rect 65616 17274 65668 17280
rect 65720 16574 65748 18022
rect 65628 16546 65748 16574
rect 65628 15570 65656 16546
rect 65616 15564 65668 15570
rect 65616 15506 65668 15512
rect 65524 14612 65576 14618
rect 65524 14554 65576 14560
rect 65628 14498 65656 15506
rect 65708 15360 65760 15366
rect 65708 15302 65760 15308
rect 65536 14470 65656 14498
rect 65536 13394 65564 14470
rect 65616 14408 65668 14414
rect 65616 14350 65668 14356
rect 65524 13388 65576 13394
rect 65524 13330 65576 13336
rect 65524 12776 65576 12782
rect 65524 12718 65576 12724
rect 65536 11642 65564 12718
rect 65628 11898 65656 14350
rect 65616 11892 65668 11898
rect 65616 11834 65668 11840
rect 65536 11614 65656 11642
rect 65524 11552 65576 11558
rect 65524 11494 65576 11500
rect 65536 3738 65564 11494
rect 65628 10606 65656 11614
rect 65616 10600 65668 10606
rect 65616 10542 65668 10548
rect 65616 10464 65668 10470
rect 65616 10406 65668 10412
rect 65524 3732 65576 3738
rect 65524 3674 65576 3680
rect 65432 876 65484 882
rect 65432 818 65484 824
rect 65248 672 65300 678
rect 65248 614 65300 620
rect 64972 604 65024 610
rect 64972 546 65024 552
rect 65338 0 65394 800
rect 65628 338 65656 10406
rect 65720 4826 65748 15302
rect 65812 7478 65840 27406
rect 65800 7472 65852 7478
rect 65800 7414 65852 7420
rect 65800 6384 65852 6390
rect 65798 6352 65800 6361
rect 65852 6352 65854 6361
rect 65798 6287 65854 6296
rect 65708 4820 65760 4826
rect 65708 4762 65760 4768
rect 65904 1358 65932 74054
rect 65984 65680 66036 65686
rect 65984 65622 66036 65628
rect 65996 50522 66024 65622
rect 66076 65408 66128 65414
rect 66076 65350 66128 65356
rect 65984 50516 66036 50522
rect 65984 50458 66036 50464
rect 65984 43784 66036 43790
rect 65984 43726 66036 43732
rect 65996 40390 66024 43726
rect 65984 40384 66036 40390
rect 65984 40326 66036 40332
rect 65982 40216 66038 40225
rect 65982 40151 66038 40160
rect 65996 38486 66024 40151
rect 65984 38480 66036 38486
rect 65984 38422 66036 38428
rect 65984 36168 66036 36174
rect 65984 36110 66036 36116
rect 65996 28218 66024 36110
rect 65984 28212 66036 28218
rect 65984 28154 66036 28160
rect 65984 25288 66036 25294
rect 65984 25230 66036 25236
rect 65996 20058 66024 25230
rect 65984 20052 66036 20058
rect 65984 19994 66036 20000
rect 65984 19916 66036 19922
rect 65984 19858 66036 19864
rect 65892 1352 65944 1358
rect 65892 1294 65944 1300
rect 65800 1284 65852 1290
rect 65800 1226 65852 1232
rect 65812 800 65840 1226
rect 65996 1018 66024 19858
rect 66088 7342 66116 65350
rect 68008 63368 68060 63374
rect 68008 63310 68060 63316
rect 66536 61736 66588 61742
rect 66536 61678 66588 61684
rect 66168 61328 66220 61334
rect 66168 61270 66220 61276
rect 66180 47258 66208 61270
rect 66260 58472 66312 58478
rect 66260 58414 66312 58420
rect 66168 47252 66220 47258
rect 66168 47194 66220 47200
rect 66168 42832 66220 42838
rect 66168 42774 66220 42780
rect 66180 33114 66208 42774
rect 66272 39642 66300 58414
rect 66352 53032 66404 53038
rect 66352 52974 66404 52980
rect 66260 39636 66312 39642
rect 66260 39578 66312 39584
rect 66260 38480 66312 38486
rect 66260 38422 66312 38428
rect 66272 34202 66300 38422
rect 66364 36378 66392 52974
rect 66444 43852 66496 43858
rect 66444 43794 66496 43800
rect 66352 36372 66404 36378
rect 66352 36314 66404 36320
rect 66352 34536 66404 34542
rect 66352 34478 66404 34484
rect 66260 34196 66312 34202
rect 66260 34138 66312 34144
rect 66168 33108 66220 33114
rect 66168 33050 66220 33056
rect 66260 30048 66312 30054
rect 66260 29990 66312 29996
rect 66168 29640 66220 29646
rect 66168 29582 66220 29588
rect 66180 16250 66208 29582
rect 66272 29306 66300 29990
rect 66260 29300 66312 29306
rect 66260 29242 66312 29248
rect 66364 29186 66392 34478
rect 66456 29850 66484 43794
rect 66548 41818 66576 61678
rect 67088 60104 67140 60110
rect 67088 60046 67140 60052
rect 66628 46980 66680 46986
rect 66628 46922 66680 46928
rect 66640 44198 66668 46922
rect 66996 45620 67048 45626
rect 66996 45562 67048 45568
rect 66812 44872 66864 44878
rect 66812 44814 66864 44820
rect 66628 44192 66680 44198
rect 66628 44134 66680 44140
rect 66720 42152 66772 42158
rect 66720 42094 66772 42100
rect 66536 41812 66588 41818
rect 66536 41754 66588 41760
rect 66536 40520 66588 40526
rect 66536 40462 66588 40468
rect 66444 29844 66496 29850
rect 66444 29786 66496 29792
rect 66444 29572 66496 29578
rect 66444 29514 66496 29520
rect 66272 29158 66392 29186
rect 66272 24886 66300 29158
rect 66352 29096 66404 29102
rect 66352 29038 66404 29044
rect 66260 24880 66312 24886
rect 66260 24822 66312 24828
rect 66364 24818 66392 29038
rect 66456 26874 66484 29514
rect 66548 27062 66576 40462
rect 66628 39976 66680 39982
rect 66628 39918 66680 39924
rect 66640 29866 66668 39918
rect 66732 30054 66760 42094
rect 66824 34746 66852 44814
rect 66904 36712 66956 36718
rect 66904 36654 66956 36660
rect 66812 34740 66864 34746
rect 66812 34682 66864 34688
rect 66812 34536 66864 34542
rect 66812 34478 66864 34484
rect 66720 30048 66772 30054
rect 66720 29990 66772 29996
rect 66640 29838 66760 29866
rect 66628 28484 66680 28490
rect 66628 28426 66680 28432
rect 66640 27878 66668 28426
rect 66628 27872 66680 27878
rect 66628 27814 66680 27820
rect 66732 27606 66760 29838
rect 66720 27600 66772 27606
rect 66720 27542 66772 27548
rect 66536 27056 66588 27062
rect 66536 26998 66588 27004
rect 66456 26846 66576 26874
rect 66444 26784 66496 26790
rect 66444 26726 66496 26732
rect 66352 24812 66404 24818
rect 66352 24754 66404 24760
rect 66260 24744 66312 24750
rect 66260 24686 66312 24692
rect 66272 20806 66300 24686
rect 66352 24200 66404 24206
rect 66352 24142 66404 24148
rect 66260 20800 66312 20806
rect 66260 20742 66312 20748
rect 66260 17128 66312 17134
rect 66260 17070 66312 17076
rect 66168 16244 66220 16250
rect 66168 16186 66220 16192
rect 66272 15366 66300 17070
rect 66260 15360 66312 15366
rect 66260 15302 66312 15308
rect 66168 12640 66220 12646
rect 66168 12582 66220 12588
rect 66076 7336 66128 7342
rect 66076 7278 66128 7284
rect 66180 5574 66208 12582
rect 66364 7818 66392 24142
rect 66456 22098 66484 26726
rect 66548 26234 66576 26846
rect 66548 26206 66760 26234
rect 66536 24268 66588 24274
rect 66536 24210 66588 24216
rect 66444 22092 66496 22098
rect 66444 22034 66496 22040
rect 66548 20346 66576 24210
rect 66628 23656 66680 23662
rect 66628 23598 66680 23604
rect 66456 20318 66576 20346
rect 66352 7812 66404 7818
rect 66352 7754 66404 7760
rect 66168 5568 66220 5574
rect 66168 5510 66220 5516
rect 66456 4758 66484 20318
rect 66640 20074 66668 23598
rect 66732 23322 66760 26206
rect 66824 23866 66852 34478
rect 66916 24410 66944 36654
rect 67008 35834 67036 45562
rect 67100 40730 67128 60046
rect 67548 51944 67600 51950
rect 67548 51886 67600 51892
rect 67560 51074 67588 51886
rect 67560 51046 67956 51074
rect 67640 50380 67692 50386
rect 67640 50322 67692 50328
rect 67180 45416 67232 45422
rect 67180 45358 67232 45364
rect 67088 40724 67140 40730
rect 67088 40666 67140 40672
rect 66996 35828 67048 35834
rect 66996 35770 67048 35776
rect 67088 34060 67140 34066
rect 67088 34002 67140 34008
rect 66996 33992 67048 33998
rect 66996 33934 67048 33940
rect 66904 24404 66956 24410
rect 66904 24346 66956 24352
rect 66812 23860 66864 23866
rect 66812 23802 66864 23808
rect 66812 23656 66864 23662
rect 66812 23598 66864 23604
rect 66720 23316 66772 23322
rect 66720 23258 66772 23264
rect 66720 22568 66772 22574
rect 66720 22510 66772 22516
rect 66548 20046 66668 20074
rect 66444 4752 66496 4758
rect 66444 4694 66496 4700
rect 66548 4554 66576 20046
rect 66628 19984 66680 19990
rect 66628 19926 66680 19932
rect 66640 5681 66668 19926
rect 66732 6730 66760 22510
rect 66824 8022 66852 23598
rect 67008 23254 67036 33934
rect 67100 25430 67128 34002
rect 67192 30938 67220 45358
rect 67272 45280 67324 45286
rect 67272 45222 67324 45228
rect 67284 34678 67312 45222
rect 67548 39432 67600 39438
rect 67548 39374 67600 39380
rect 67456 37256 67508 37262
rect 67456 37198 67508 37204
rect 67364 36236 67416 36242
rect 67364 36178 67416 36184
rect 67272 34672 67324 34678
rect 67272 34614 67324 34620
rect 67272 31952 67324 31958
rect 67272 31894 67324 31900
rect 67180 30932 67232 30938
rect 67180 30874 67232 30880
rect 67180 30184 67232 30190
rect 67180 30126 67232 30132
rect 67088 25424 67140 25430
rect 67088 25366 67140 25372
rect 67088 25288 67140 25294
rect 67088 25230 67140 25236
rect 66996 23248 67048 23254
rect 66996 23190 67048 23196
rect 66904 23112 66956 23118
rect 66904 23054 66956 23060
rect 66812 8016 66864 8022
rect 66812 7958 66864 7964
rect 66916 6798 66944 23054
rect 66996 20324 67048 20330
rect 66996 20266 67048 20272
rect 67008 16114 67036 20266
rect 67100 19990 67128 25230
rect 67088 19984 67140 19990
rect 67088 19926 67140 19932
rect 66996 16108 67048 16114
rect 66996 16050 67048 16056
rect 67192 7546 67220 30126
rect 67284 29102 67312 31894
rect 67272 29096 67324 29102
rect 67272 29038 67324 29044
rect 67272 28960 67324 28966
rect 67272 28902 67324 28908
rect 67284 27130 67312 28902
rect 67272 27124 67324 27130
rect 67272 27066 67324 27072
rect 67272 26376 67324 26382
rect 67272 26318 67324 26324
rect 67180 7540 67232 7546
rect 67180 7482 67232 7488
rect 66904 6792 66956 6798
rect 66904 6734 66956 6740
rect 66720 6724 66772 6730
rect 66720 6666 66772 6672
rect 66626 5672 66682 5681
rect 66626 5607 66682 5616
rect 67284 4690 67312 26318
rect 67376 24682 67404 36178
rect 67468 25498 67496 37198
rect 67456 25492 67508 25498
rect 67456 25434 67508 25440
rect 67456 25356 67508 25362
rect 67456 25298 67508 25304
rect 67364 24676 67416 24682
rect 67364 24618 67416 24624
rect 67364 23180 67416 23186
rect 67364 23122 67416 23128
rect 67376 6322 67404 23122
rect 67468 23050 67496 25298
rect 67456 23044 67508 23050
rect 67456 22986 67508 22992
rect 67456 20800 67508 20806
rect 67456 20742 67508 20748
rect 67468 7410 67496 20742
rect 67560 20602 67588 39374
rect 67652 34202 67680 50322
rect 67928 35290 67956 51046
rect 68020 42770 68048 63310
rect 68008 42764 68060 42770
rect 68008 42706 68060 42712
rect 67916 35284 67968 35290
rect 67916 35226 67968 35232
rect 67732 34536 67784 34542
rect 67732 34478 67784 34484
rect 67640 34196 67692 34202
rect 67640 34138 67692 34144
rect 67744 23866 67772 34478
rect 67824 31816 67876 31822
rect 67824 31758 67876 31764
rect 67732 23860 67784 23866
rect 67732 23802 67784 23808
rect 67640 22024 67692 22030
rect 67640 21966 67692 21972
rect 67548 20596 67600 20602
rect 67548 20538 67600 20544
rect 67548 15360 67600 15366
rect 67548 15302 67600 15308
rect 67560 8090 67588 15302
rect 67548 8084 67600 8090
rect 67548 8026 67600 8032
rect 67456 7404 67508 7410
rect 67456 7346 67508 7352
rect 67364 6316 67416 6322
rect 67364 6258 67416 6264
rect 67652 5710 67680 21966
rect 67836 16590 67864 31758
rect 68008 28008 68060 28014
rect 68008 27950 68060 27956
rect 67916 23112 67968 23118
rect 67916 23054 67968 23060
rect 67824 16584 67876 16590
rect 67824 16526 67876 16532
rect 67732 14408 67784 14414
rect 67732 14350 67784 14356
rect 67640 5704 67692 5710
rect 67640 5646 67692 5652
rect 67744 5370 67772 14350
rect 67928 7002 67956 23054
rect 67916 6996 67968 7002
rect 67916 6938 67968 6944
rect 68020 6458 68048 27950
rect 68112 16574 68140 76434
rect 68560 41608 68612 41614
rect 68560 41550 68612 41556
rect 68192 40520 68244 40526
rect 68192 40462 68244 40468
rect 68204 21146 68232 40462
rect 68284 36168 68336 36174
rect 68284 36110 68336 36116
rect 68192 21140 68244 21146
rect 68192 21082 68244 21088
rect 68296 20618 68324 36110
rect 68376 35624 68428 35630
rect 68376 35566 68428 35572
rect 68388 24410 68416 35566
rect 68468 35080 68520 35086
rect 68468 35022 68520 35028
rect 68376 24404 68428 24410
rect 68376 24346 68428 24352
rect 68204 20590 68324 20618
rect 68204 19514 68232 20590
rect 68284 20460 68336 20466
rect 68284 20402 68336 20408
rect 68192 19508 68244 19514
rect 68192 19450 68244 19456
rect 68112 16546 68232 16574
rect 68100 13320 68152 13326
rect 68100 13262 68152 13268
rect 68008 6452 68060 6458
rect 68008 6394 68060 6400
rect 67732 5364 67784 5370
rect 67732 5306 67784 5312
rect 67272 4684 67324 4690
rect 67272 4626 67324 4632
rect 66536 4548 66588 4554
rect 66536 4490 66588 4496
rect 68112 4214 68140 13262
rect 68100 4208 68152 4214
rect 68100 4150 68152 4156
rect 66812 3052 66864 3058
rect 66812 2994 66864 3000
rect 66260 2848 66312 2854
rect 66260 2790 66312 2796
rect 66272 2650 66300 2790
rect 66260 2644 66312 2650
rect 66260 2586 66312 2592
rect 66076 2440 66128 2446
rect 66076 2382 66128 2388
rect 66088 2106 66116 2382
rect 66076 2100 66128 2106
rect 66076 2042 66128 2048
rect 66824 1970 66852 2994
rect 66996 2848 67048 2854
rect 66996 2790 67048 2796
rect 67008 2514 67036 2790
rect 66996 2508 67048 2514
rect 66996 2450 67048 2456
rect 67088 2440 67140 2446
rect 67088 2382 67140 2388
rect 66812 1964 66864 1970
rect 66812 1906 66864 1912
rect 65984 1012 66036 1018
rect 65984 954 66036 960
rect 66732 870 66852 898
rect 66732 800 66760 870
rect 65616 332 65668 338
rect 65616 274 65668 280
rect 65798 0 65854 800
rect 66258 0 66314 800
rect 66718 0 66774 800
rect 66824 762 66852 870
rect 67100 762 67128 2382
rect 68100 2304 68152 2310
rect 68100 2246 68152 2252
rect 68112 1970 68140 2246
rect 68100 1964 68152 1970
rect 68100 1906 68152 1912
rect 67456 1760 67508 1766
rect 67456 1702 67508 1708
rect 67180 1420 67232 1426
rect 67180 1362 67232 1368
rect 67192 800 67220 1362
rect 67468 1358 67496 1702
rect 68204 1358 68232 16546
rect 68296 2038 68324 20402
rect 68376 20392 68428 20398
rect 68376 20334 68428 20340
rect 68388 3126 68416 20334
rect 68480 18970 68508 35022
rect 68572 22098 68600 41550
rect 68560 22092 68612 22098
rect 68560 22034 68612 22040
rect 68560 19304 68612 19310
rect 68560 19246 68612 19252
rect 68468 18964 68520 18970
rect 68468 18906 68520 18912
rect 68376 3120 68428 3126
rect 68376 3062 68428 3068
rect 68468 2848 68520 2854
rect 68468 2790 68520 2796
rect 68480 2514 68508 2790
rect 68468 2508 68520 2514
rect 68468 2450 68520 2456
rect 68376 2440 68428 2446
rect 68376 2382 68428 2388
rect 68284 2032 68336 2038
rect 68284 1974 68336 1980
rect 67456 1352 67508 1358
rect 67456 1294 67508 1300
rect 68192 1352 68244 1358
rect 68192 1294 68244 1300
rect 68112 870 68232 898
rect 68112 800 68140 870
rect 66824 734 67128 762
rect 67178 0 67234 800
rect 67638 0 67694 800
rect 68098 0 68154 800
rect 68204 762 68232 870
rect 68388 762 68416 2382
rect 68572 1986 68600 19246
rect 68480 1958 68600 1986
rect 68664 1970 68692 78610
rect 69296 56840 69348 56846
rect 69296 56782 69348 56788
rect 69112 55276 69164 55282
rect 69112 55218 69164 55224
rect 69020 53440 69072 53446
rect 69020 53382 69072 53388
rect 69032 35154 69060 53382
rect 69124 38010 69152 55218
rect 69204 48136 69256 48142
rect 69204 48078 69256 48084
rect 69112 38004 69164 38010
rect 69112 37946 69164 37952
rect 69020 35148 69072 35154
rect 69020 35090 69072 35096
rect 68836 33992 68888 33998
rect 68836 33934 68888 33940
rect 68744 26920 68796 26926
rect 68744 26862 68796 26868
rect 68756 7206 68784 26862
rect 68848 17882 68876 33934
rect 69112 28756 69164 28762
rect 69112 28698 69164 28704
rect 69020 27872 69072 27878
rect 69020 27814 69072 27820
rect 68928 23656 68980 23662
rect 68928 23598 68980 23604
rect 68836 17876 68888 17882
rect 68836 17818 68888 17824
rect 68744 7200 68796 7206
rect 68744 7142 68796 7148
rect 68940 6662 68968 23598
rect 68928 6656 68980 6662
rect 68928 6598 68980 6604
rect 69032 3369 69060 27814
rect 69124 5234 69152 28698
rect 69216 26586 69244 48078
rect 69308 38554 69336 56782
rect 69388 53576 69440 53582
rect 69388 53518 69440 53524
rect 69296 38548 69348 38554
rect 69296 38490 69348 38496
rect 69400 35766 69428 53518
rect 69756 48816 69808 48822
rect 69756 48758 69808 48764
rect 69572 48680 69624 48686
rect 69572 48622 69624 48628
rect 69480 38344 69532 38350
rect 69480 38286 69532 38292
rect 69388 35760 69440 35766
rect 69388 35702 69440 35708
rect 69296 32904 69348 32910
rect 69296 32846 69348 32852
rect 69204 26580 69256 26586
rect 69204 26522 69256 26528
rect 69204 18216 69256 18222
rect 69204 18158 69256 18164
rect 69216 11778 69244 18158
rect 69308 11914 69336 32846
rect 69388 31272 69440 31278
rect 69388 31214 69440 31220
rect 69400 14550 69428 31214
rect 69492 20534 69520 38286
rect 69584 32570 69612 48622
rect 69664 47048 69716 47054
rect 69664 46990 69716 46996
rect 69572 32564 69624 32570
rect 69572 32506 69624 32512
rect 69676 32026 69704 46990
rect 69664 32020 69716 32026
rect 69664 31962 69716 31968
rect 69664 30728 69716 30734
rect 69664 30670 69716 30676
rect 69572 29164 69624 29170
rect 69572 29106 69624 29112
rect 69480 20528 69532 20534
rect 69480 20470 69532 20476
rect 69480 19848 69532 19854
rect 69480 19790 69532 19796
rect 69388 14544 69440 14550
rect 69388 14486 69440 14492
rect 69492 12322 69520 19790
rect 69584 15162 69612 29106
rect 69676 15706 69704 30670
rect 69768 27402 69796 48758
rect 70124 42696 70176 42702
rect 70124 42638 70176 42644
rect 69848 38888 69900 38894
rect 69848 38830 69900 38836
rect 69756 27396 69808 27402
rect 69756 27338 69808 27344
rect 69860 26042 69888 38830
rect 70032 37800 70084 37806
rect 70032 37742 70084 37748
rect 69848 26036 69900 26042
rect 69848 25978 69900 25984
rect 69756 24744 69808 24750
rect 69756 24686 69808 24692
rect 69664 15700 69716 15706
rect 69664 15642 69716 15648
rect 69572 15156 69624 15162
rect 69572 15098 69624 15104
rect 69664 14952 69716 14958
rect 69664 14894 69716 14900
rect 69572 14544 69624 14550
rect 69572 14486 69624 14492
rect 69400 12294 69520 12322
rect 69400 12050 69428 12294
rect 69400 12022 69520 12050
rect 69308 11886 69428 11914
rect 69216 11750 69336 11778
rect 69204 11688 69256 11694
rect 69204 11630 69256 11636
rect 69216 6118 69244 11630
rect 69204 6112 69256 6118
rect 69204 6054 69256 6060
rect 69308 5302 69336 11750
rect 69296 5296 69348 5302
rect 69296 5238 69348 5244
rect 69112 5228 69164 5234
rect 69112 5170 69164 5176
rect 69400 5098 69428 11886
rect 69492 5642 69520 12022
rect 69480 5636 69532 5642
rect 69480 5578 69532 5584
rect 69584 5166 69612 14486
rect 69572 5160 69624 5166
rect 69572 5102 69624 5108
rect 69388 5092 69440 5098
rect 69388 5034 69440 5040
rect 69018 3360 69074 3369
rect 69018 3295 69074 3304
rect 69112 3052 69164 3058
rect 69112 2994 69164 3000
rect 69020 2984 69072 2990
rect 69020 2926 69072 2932
rect 69032 2106 69060 2926
rect 69124 2650 69152 2994
rect 69480 2984 69532 2990
rect 69480 2926 69532 2932
rect 69388 2916 69440 2922
rect 69388 2858 69440 2864
rect 69112 2644 69164 2650
rect 69112 2586 69164 2592
rect 69020 2100 69072 2106
rect 69020 2042 69072 2048
rect 68652 1964 68704 1970
rect 68480 1562 68508 1958
rect 68652 1906 68704 1912
rect 68560 1896 68612 1902
rect 68560 1838 68612 1844
rect 68468 1556 68520 1562
rect 68468 1498 68520 1504
rect 68572 800 68600 1838
rect 69400 1358 69428 2858
rect 69388 1352 69440 1358
rect 69388 1294 69440 1300
rect 69492 800 69520 2926
rect 69676 2582 69704 14894
rect 69768 5778 69796 24686
rect 69940 22024 69992 22030
rect 69940 21966 69992 21972
rect 69848 21480 69900 21486
rect 69848 21422 69900 21428
rect 69860 6390 69888 21422
rect 69848 6384 69900 6390
rect 69848 6326 69900 6332
rect 69756 5772 69808 5778
rect 69756 5714 69808 5720
rect 69952 5574 69980 21966
rect 70044 20262 70072 37742
rect 70136 22098 70164 42638
rect 70216 32360 70268 32366
rect 70216 32302 70268 32308
rect 70124 22092 70176 22098
rect 70124 22034 70176 22040
rect 70124 20936 70176 20942
rect 70124 20878 70176 20884
rect 70032 20256 70084 20262
rect 70032 20198 70084 20204
rect 69940 5568 69992 5574
rect 69940 5510 69992 5516
rect 69664 2576 69716 2582
rect 69664 2518 69716 2524
rect 70136 2514 70164 20878
rect 70228 17338 70256 32302
rect 70584 17672 70636 17678
rect 70584 17614 70636 17620
rect 70216 17332 70268 17338
rect 70216 17274 70268 17280
rect 70492 17196 70544 17202
rect 70492 17138 70544 17144
rect 70400 16040 70452 16046
rect 70400 15982 70452 15988
rect 70412 6866 70440 15982
rect 70400 6860 70452 6866
rect 70400 6802 70452 6808
rect 70124 2508 70176 2514
rect 70124 2450 70176 2456
rect 69756 2304 69808 2310
rect 69756 2246 69808 2252
rect 69768 1358 69796 2246
rect 69940 1420 69992 1426
rect 69940 1362 69992 1368
rect 69756 1352 69808 1358
rect 69756 1294 69808 1300
rect 69952 800 69980 1362
rect 68204 734 68416 762
rect 68558 0 68614 800
rect 69018 0 69074 800
rect 69478 0 69534 800
rect 69938 0 69994 800
rect 70398 0 70454 800
rect 70504 746 70532 17138
rect 70596 3466 70624 17614
rect 70688 6914 70716 80786
rect 71136 69964 71188 69970
rect 71136 69906 71188 69912
rect 70768 47116 70820 47122
rect 70768 47058 70820 47064
rect 70780 15366 70808 47058
rect 70860 44192 70912 44198
rect 70860 44134 70912 44140
rect 70768 15360 70820 15366
rect 70768 15302 70820 15308
rect 70872 11150 70900 44134
rect 70952 15496 71004 15502
rect 70952 15438 71004 15444
rect 70860 11144 70912 11150
rect 70860 11086 70912 11092
rect 70688 6886 70808 6914
rect 70584 3460 70636 3466
rect 70584 3402 70636 3408
rect 70676 2916 70728 2922
rect 70676 2858 70728 2864
rect 70688 2514 70716 2858
rect 70676 2508 70728 2514
rect 70676 2450 70728 2456
rect 70676 2304 70728 2310
rect 70676 2246 70728 2252
rect 70688 1970 70716 2246
rect 70676 1964 70728 1970
rect 70676 1906 70728 1912
rect 70780 1358 70808 6886
rect 70964 3194 70992 15438
rect 71148 6914 71176 69906
rect 71320 59084 71372 59090
rect 71320 59026 71372 59032
rect 71228 54664 71280 54670
rect 71228 54606 71280 54612
rect 71056 6886 71176 6914
rect 70952 3188 71004 3194
rect 70952 3130 71004 3136
rect 71056 3074 71084 6886
rect 71136 5568 71188 5574
rect 71136 5510 71188 5516
rect 70964 3046 71084 3074
rect 70860 2848 70912 2854
rect 70860 2790 70912 2796
rect 70872 1970 70900 2790
rect 70860 1964 70912 1970
rect 70860 1906 70912 1912
rect 70964 1834 70992 3046
rect 71044 2984 71096 2990
rect 71044 2926 71096 2932
rect 71056 2650 71084 2926
rect 71044 2644 71096 2650
rect 71044 2586 71096 2592
rect 71148 2038 71176 5510
rect 71240 2582 71268 54606
rect 71332 6225 71360 59026
rect 71504 25832 71556 25838
rect 71504 25774 71556 25780
rect 71318 6216 71374 6225
rect 71318 6151 71374 6160
rect 71516 5846 71544 25774
rect 71596 22024 71648 22030
rect 71596 21966 71648 21972
rect 71504 5840 71556 5846
rect 71504 5782 71556 5788
rect 71608 5574 71636 21966
rect 71596 5568 71648 5574
rect 71596 5510 71648 5516
rect 71228 2576 71280 2582
rect 71228 2518 71280 2524
rect 71136 2032 71188 2038
rect 71136 1974 71188 1980
rect 71700 1970 71728 82962
rect 71836 82236 72188 83206
rect 71836 82180 71864 82236
rect 71920 82180 71944 82236
rect 72000 82180 72024 82236
rect 72080 82180 72104 82236
rect 72160 82180 72188 82236
rect 71836 82170 72188 82180
rect 71836 82118 71858 82170
rect 71910 82156 71922 82170
rect 71974 82156 71986 82170
rect 72038 82156 72050 82170
rect 72102 82156 72114 82170
rect 71920 82118 71922 82156
rect 72102 82118 72104 82156
rect 72166 82118 72188 82170
rect 71836 82100 71864 82118
rect 71920 82100 71944 82118
rect 72000 82100 72024 82118
rect 72080 82100 72104 82118
rect 72160 82100 72188 82118
rect 71836 82076 72188 82100
rect 71836 82020 71864 82076
rect 71920 82020 71944 82076
rect 72000 82020 72024 82076
rect 72080 82020 72104 82076
rect 72160 82020 72188 82076
rect 71836 81996 72188 82020
rect 71836 81940 71864 81996
rect 71920 81940 71944 81996
rect 72000 81940 72024 81996
rect 72080 81940 72104 81996
rect 72160 81940 72188 81996
rect 71836 81082 72188 81940
rect 71836 81030 71858 81082
rect 71910 81030 71922 81082
rect 71974 81030 71986 81082
rect 72038 81030 72050 81082
rect 72102 81030 72114 81082
rect 72166 81030 72188 81082
rect 71836 79994 72188 81030
rect 71836 79942 71858 79994
rect 71910 79942 71922 79994
rect 71974 79942 71986 79994
rect 72038 79942 72050 79994
rect 72102 79942 72114 79994
rect 72166 79942 72188 79994
rect 71836 78906 72188 79942
rect 71836 78854 71858 78906
rect 71910 78854 71922 78906
rect 71974 78854 71986 78906
rect 72038 78854 72050 78906
rect 72102 78854 72114 78906
rect 72166 78854 72188 78906
rect 71836 77818 72188 78854
rect 71836 77766 71858 77818
rect 71910 77766 71922 77818
rect 71974 77766 71986 77818
rect 72038 77766 72050 77818
rect 72102 77766 72114 77818
rect 72166 77766 72188 77818
rect 71836 76730 72188 77766
rect 71836 76678 71858 76730
rect 71910 76678 71922 76730
rect 71974 76678 71986 76730
rect 72038 76678 72050 76730
rect 72102 76678 72114 76730
rect 72166 76678 72188 76730
rect 71836 75642 72188 76678
rect 71836 75590 71858 75642
rect 71910 75590 71922 75642
rect 71974 75590 71986 75642
rect 72038 75590 72050 75642
rect 72102 75590 72114 75642
rect 72166 75590 72188 75642
rect 71836 74554 72188 75590
rect 71836 74502 71858 74554
rect 71910 74502 71922 74554
rect 71974 74502 71986 74554
rect 72038 74502 72050 74554
rect 72102 74502 72114 74554
rect 72166 74502 72188 74554
rect 71836 73466 72188 74502
rect 71836 73414 71858 73466
rect 71910 73414 71922 73466
rect 71974 73414 71986 73466
rect 72038 73414 72050 73466
rect 72102 73414 72114 73466
rect 72166 73414 72188 73466
rect 71836 72378 72188 73414
rect 71836 72326 71858 72378
rect 71910 72326 71922 72378
rect 71974 72326 71986 72378
rect 72038 72326 72050 72378
rect 72102 72326 72114 72378
rect 72166 72326 72188 72378
rect 71836 72236 72188 72326
rect 71836 72180 71864 72236
rect 71920 72180 71944 72236
rect 72000 72180 72024 72236
rect 72080 72180 72104 72236
rect 72160 72180 72188 72236
rect 71836 72156 72188 72180
rect 71836 72100 71864 72156
rect 71920 72100 71944 72156
rect 72000 72100 72024 72156
rect 72080 72100 72104 72156
rect 72160 72100 72188 72156
rect 71836 72076 72188 72100
rect 71836 72020 71864 72076
rect 71920 72020 71944 72076
rect 72000 72020 72024 72076
rect 72080 72020 72104 72076
rect 72160 72020 72188 72076
rect 71836 71996 72188 72020
rect 71836 71940 71864 71996
rect 71920 71940 71944 71996
rect 72000 71940 72024 71996
rect 72080 71940 72104 71996
rect 72160 71940 72188 71996
rect 71836 71290 72188 71940
rect 71836 71238 71858 71290
rect 71910 71238 71922 71290
rect 71974 71238 71986 71290
rect 72038 71238 72050 71290
rect 72102 71238 72114 71290
rect 72166 71238 72188 71290
rect 71836 70202 72188 71238
rect 71836 70150 71858 70202
rect 71910 70150 71922 70202
rect 71974 70150 71986 70202
rect 72038 70150 72050 70202
rect 72102 70150 72114 70202
rect 72166 70150 72188 70202
rect 71836 69114 72188 70150
rect 71836 69062 71858 69114
rect 71910 69062 71922 69114
rect 71974 69062 71986 69114
rect 72038 69062 72050 69114
rect 72102 69062 72114 69114
rect 72166 69062 72188 69114
rect 71836 68026 72188 69062
rect 71836 67974 71858 68026
rect 71910 67974 71922 68026
rect 71974 67974 71986 68026
rect 72038 67974 72050 68026
rect 72102 67974 72114 68026
rect 72166 67974 72188 68026
rect 71836 66938 72188 67974
rect 74188 85978 74540 86000
rect 74188 85926 74210 85978
rect 74262 85926 74274 85978
rect 74326 85926 74338 85978
rect 74390 85926 74402 85978
rect 74454 85926 74466 85978
rect 74518 85926 74540 85978
rect 74188 84890 74540 85926
rect 74188 84838 74210 84890
rect 74262 84838 74274 84890
rect 74326 84838 74338 84890
rect 74390 84838 74402 84890
rect 74454 84838 74466 84890
rect 74518 84838 74540 84890
rect 74188 84588 74540 84838
rect 74188 84532 74216 84588
rect 74272 84532 74296 84588
rect 74352 84532 74376 84588
rect 74432 84532 74456 84588
rect 74512 84532 74540 84588
rect 74188 84508 74540 84532
rect 74188 84452 74216 84508
rect 74272 84452 74296 84508
rect 74352 84452 74376 84508
rect 74432 84452 74456 84508
rect 74512 84452 74540 84508
rect 74188 84428 74540 84452
rect 74188 84372 74216 84428
rect 74272 84372 74296 84428
rect 74352 84372 74376 84428
rect 74432 84372 74456 84428
rect 74512 84372 74540 84428
rect 74188 84348 74540 84372
rect 74188 84292 74216 84348
rect 74272 84292 74296 84348
rect 74352 84292 74376 84348
rect 74432 84292 74456 84348
rect 74512 84292 74540 84348
rect 74188 83802 74540 84292
rect 74188 83750 74210 83802
rect 74262 83750 74274 83802
rect 74326 83750 74338 83802
rect 74390 83750 74402 83802
rect 74454 83750 74466 83802
rect 74518 83750 74540 83802
rect 74188 82714 74540 83750
rect 74188 82662 74210 82714
rect 74262 82662 74274 82714
rect 74326 82662 74338 82714
rect 74390 82662 74402 82714
rect 74454 82662 74466 82714
rect 74518 82662 74540 82714
rect 74188 81626 74540 82662
rect 74188 81574 74210 81626
rect 74262 81574 74274 81626
rect 74326 81574 74338 81626
rect 74390 81574 74402 81626
rect 74454 81574 74466 81626
rect 74518 81574 74540 81626
rect 74188 80538 74540 81574
rect 74188 80486 74210 80538
rect 74262 80486 74274 80538
rect 74326 80486 74338 80538
rect 74390 80486 74402 80538
rect 74454 80486 74466 80538
rect 74518 80486 74540 80538
rect 74188 79450 74540 80486
rect 74188 79398 74210 79450
rect 74262 79398 74274 79450
rect 74326 79398 74338 79450
rect 74390 79398 74402 79450
rect 74454 79398 74466 79450
rect 74518 79398 74540 79450
rect 74188 78362 74540 79398
rect 74188 78310 74210 78362
rect 74262 78310 74274 78362
rect 74326 78310 74338 78362
rect 74390 78310 74402 78362
rect 74454 78310 74466 78362
rect 74518 78310 74540 78362
rect 74188 77274 74540 78310
rect 74188 77222 74210 77274
rect 74262 77222 74274 77274
rect 74326 77222 74338 77274
rect 74390 77222 74402 77274
rect 74454 77222 74466 77274
rect 74518 77222 74540 77274
rect 74188 76186 74540 77222
rect 74188 76134 74210 76186
rect 74262 76134 74274 76186
rect 74326 76134 74338 76186
rect 74390 76134 74402 76186
rect 74454 76134 74466 76186
rect 74518 76134 74540 76186
rect 74188 75098 74540 76134
rect 74188 75046 74210 75098
rect 74262 75046 74274 75098
rect 74326 75046 74338 75098
rect 74390 75046 74402 75098
rect 74454 75046 74466 75098
rect 74518 75046 74540 75098
rect 74188 74588 74540 75046
rect 74188 74532 74216 74588
rect 74272 74532 74296 74588
rect 74352 74532 74376 74588
rect 74432 74532 74456 74588
rect 74512 74532 74540 74588
rect 74188 74508 74540 74532
rect 74188 74452 74216 74508
rect 74272 74452 74296 74508
rect 74352 74452 74376 74508
rect 74432 74452 74456 74508
rect 74512 74452 74540 74508
rect 74188 74428 74540 74452
rect 74188 74372 74216 74428
rect 74272 74372 74296 74428
rect 74352 74372 74376 74428
rect 74432 74372 74456 74428
rect 74512 74372 74540 74428
rect 74188 74348 74540 74372
rect 74188 74292 74216 74348
rect 74272 74292 74296 74348
rect 74352 74292 74376 74348
rect 74432 74292 74456 74348
rect 74512 74292 74540 74348
rect 74188 74010 74540 74292
rect 74188 73958 74210 74010
rect 74262 73958 74274 74010
rect 74326 73958 74338 74010
rect 74390 73958 74402 74010
rect 74454 73958 74466 74010
rect 74518 73958 74540 74010
rect 74188 72922 74540 73958
rect 74188 72870 74210 72922
rect 74262 72870 74274 72922
rect 74326 72870 74338 72922
rect 74390 72870 74402 72922
rect 74454 72870 74466 72922
rect 74518 72870 74540 72922
rect 74188 71834 74540 72870
rect 74188 71782 74210 71834
rect 74262 71782 74274 71834
rect 74326 71782 74338 71834
rect 74390 71782 74402 71834
rect 74454 71782 74466 71834
rect 74518 71782 74540 71834
rect 74188 70746 74540 71782
rect 74188 70694 74210 70746
rect 74262 70694 74274 70746
rect 74326 70694 74338 70746
rect 74390 70694 74402 70746
rect 74454 70694 74466 70746
rect 74518 70694 74540 70746
rect 74188 69658 74540 70694
rect 74188 69606 74210 69658
rect 74262 69606 74274 69658
rect 74326 69606 74338 69658
rect 74390 69606 74402 69658
rect 74454 69606 74466 69658
rect 74518 69606 74540 69658
rect 74188 68570 74540 69606
rect 74188 68518 74210 68570
rect 74262 68518 74274 68570
rect 74326 68518 74338 68570
rect 74390 68518 74402 68570
rect 74454 68518 74466 68570
rect 74518 68518 74540 68570
rect 72792 67788 72844 67794
rect 72792 67730 72844 67736
rect 71836 66886 71858 66938
rect 71910 66886 71922 66938
rect 71974 66886 71986 66938
rect 72038 66886 72050 66938
rect 72102 66886 72114 66938
rect 72166 66886 72188 66938
rect 71836 65850 72188 66886
rect 71836 65798 71858 65850
rect 71910 65798 71922 65850
rect 71974 65798 71986 65850
rect 72038 65798 72050 65850
rect 72102 65798 72114 65850
rect 72166 65798 72188 65850
rect 71836 64762 72188 65798
rect 71836 64710 71858 64762
rect 71910 64710 71922 64762
rect 71974 64710 71986 64762
rect 72038 64710 72050 64762
rect 72102 64710 72114 64762
rect 72166 64710 72188 64762
rect 71836 63674 72188 64710
rect 71836 63622 71858 63674
rect 71910 63622 71922 63674
rect 71974 63622 71986 63674
rect 72038 63622 72050 63674
rect 72102 63622 72114 63674
rect 72166 63622 72188 63674
rect 71836 62586 72188 63622
rect 71836 62534 71858 62586
rect 71910 62534 71922 62586
rect 71974 62534 71986 62586
rect 72038 62534 72050 62586
rect 72102 62534 72114 62586
rect 72166 62534 72188 62586
rect 71836 62236 72188 62534
rect 71836 62180 71864 62236
rect 71920 62180 71944 62236
rect 72000 62180 72024 62236
rect 72080 62180 72104 62236
rect 72160 62180 72188 62236
rect 71836 62156 72188 62180
rect 71836 62100 71864 62156
rect 71920 62100 71944 62156
rect 72000 62100 72024 62156
rect 72080 62100 72104 62156
rect 72160 62100 72188 62156
rect 71836 62076 72188 62100
rect 71836 62020 71864 62076
rect 71920 62020 71944 62076
rect 72000 62020 72024 62076
rect 72080 62020 72104 62076
rect 72160 62020 72188 62076
rect 71836 61996 72188 62020
rect 71836 61940 71864 61996
rect 71920 61940 71944 61996
rect 72000 61940 72024 61996
rect 72080 61940 72104 61996
rect 72160 61940 72188 61996
rect 71836 61498 72188 61940
rect 71836 61446 71858 61498
rect 71910 61446 71922 61498
rect 71974 61446 71986 61498
rect 72038 61446 72050 61498
rect 72102 61446 72114 61498
rect 72166 61446 72188 61498
rect 71836 60410 72188 61446
rect 71836 60358 71858 60410
rect 71910 60358 71922 60410
rect 71974 60358 71986 60410
rect 72038 60358 72050 60410
rect 72102 60358 72114 60410
rect 72166 60358 72188 60410
rect 71836 59322 72188 60358
rect 71836 59270 71858 59322
rect 71910 59270 71922 59322
rect 71974 59270 71986 59322
rect 72038 59270 72050 59322
rect 72102 59270 72114 59322
rect 72166 59270 72188 59322
rect 71836 58234 72188 59270
rect 71836 58182 71858 58234
rect 71910 58182 71922 58234
rect 71974 58182 71986 58234
rect 72038 58182 72050 58234
rect 72102 58182 72114 58234
rect 72166 58182 72188 58234
rect 71836 57146 72188 58182
rect 71836 57094 71858 57146
rect 71910 57094 71922 57146
rect 71974 57094 71986 57146
rect 72038 57094 72050 57146
rect 72102 57094 72114 57146
rect 72166 57094 72188 57146
rect 71836 56058 72188 57094
rect 71836 56006 71858 56058
rect 71910 56006 71922 56058
rect 71974 56006 71986 56058
rect 72038 56006 72050 56058
rect 72102 56006 72114 56058
rect 72166 56006 72188 56058
rect 71836 54970 72188 56006
rect 71836 54918 71858 54970
rect 71910 54918 71922 54970
rect 71974 54918 71986 54970
rect 72038 54918 72050 54970
rect 72102 54918 72114 54970
rect 72166 54918 72188 54970
rect 71836 53882 72188 54918
rect 71836 53830 71858 53882
rect 71910 53830 71922 53882
rect 71974 53830 71986 53882
rect 72038 53830 72050 53882
rect 72102 53830 72114 53882
rect 72166 53830 72188 53882
rect 71836 52794 72188 53830
rect 71836 52742 71858 52794
rect 71910 52742 71922 52794
rect 71974 52742 71986 52794
rect 72038 52742 72050 52794
rect 72102 52742 72114 52794
rect 72166 52742 72188 52794
rect 71836 52236 72188 52742
rect 71836 52180 71864 52236
rect 71920 52180 71944 52236
rect 72000 52180 72024 52236
rect 72080 52180 72104 52236
rect 72160 52180 72188 52236
rect 71836 52156 72188 52180
rect 71836 52100 71864 52156
rect 71920 52100 71944 52156
rect 72000 52100 72024 52156
rect 72080 52100 72104 52156
rect 72160 52100 72188 52156
rect 71836 52076 72188 52100
rect 71836 52020 71864 52076
rect 71920 52020 71944 52076
rect 72000 52020 72024 52076
rect 72080 52020 72104 52076
rect 72160 52020 72188 52076
rect 71836 51996 72188 52020
rect 71836 51940 71864 51996
rect 71920 51940 71944 51996
rect 72000 51940 72024 51996
rect 72080 51940 72104 51996
rect 72160 51940 72188 51996
rect 71836 51706 72188 51940
rect 71836 51654 71858 51706
rect 71910 51654 71922 51706
rect 71974 51654 71986 51706
rect 72038 51654 72050 51706
rect 72102 51654 72114 51706
rect 72166 51654 72188 51706
rect 71836 50618 72188 51654
rect 71836 50566 71858 50618
rect 71910 50566 71922 50618
rect 71974 50566 71986 50618
rect 72038 50566 72050 50618
rect 72102 50566 72114 50618
rect 72166 50566 72188 50618
rect 71836 49530 72188 50566
rect 71836 49478 71858 49530
rect 71910 49478 71922 49530
rect 71974 49478 71986 49530
rect 72038 49478 72050 49530
rect 72102 49478 72114 49530
rect 72166 49478 72188 49530
rect 71836 48442 72188 49478
rect 71836 48390 71858 48442
rect 71910 48390 71922 48442
rect 71974 48390 71986 48442
rect 72038 48390 72050 48442
rect 72102 48390 72114 48442
rect 72166 48390 72188 48442
rect 71836 47354 72188 48390
rect 71836 47302 71858 47354
rect 71910 47302 71922 47354
rect 71974 47302 71986 47354
rect 72038 47302 72050 47354
rect 72102 47302 72114 47354
rect 72166 47302 72188 47354
rect 71836 46266 72188 47302
rect 71836 46214 71858 46266
rect 71910 46214 71922 46266
rect 71974 46214 71986 46266
rect 72038 46214 72050 46266
rect 72102 46214 72114 46266
rect 72166 46214 72188 46266
rect 71836 45178 72188 46214
rect 71836 45126 71858 45178
rect 71910 45126 71922 45178
rect 71974 45126 71986 45178
rect 72038 45126 72050 45178
rect 72102 45126 72114 45178
rect 72166 45126 72188 45178
rect 71836 44090 72188 45126
rect 71836 44038 71858 44090
rect 71910 44038 71922 44090
rect 71974 44038 71986 44090
rect 72038 44038 72050 44090
rect 72102 44038 72114 44090
rect 72166 44038 72188 44090
rect 71836 43002 72188 44038
rect 71836 42950 71858 43002
rect 71910 42950 71922 43002
rect 71974 42950 71986 43002
rect 72038 42950 72050 43002
rect 72102 42950 72114 43002
rect 72166 42950 72188 43002
rect 71836 42236 72188 42950
rect 71836 42180 71864 42236
rect 71920 42180 71944 42236
rect 72000 42180 72024 42236
rect 72080 42180 72104 42236
rect 72160 42180 72188 42236
rect 71836 42156 72188 42180
rect 71836 42100 71864 42156
rect 71920 42100 71944 42156
rect 72000 42100 72024 42156
rect 72080 42100 72104 42156
rect 72160 42100 72188 42156
rect 71836 42076 72188 42100
rect 71836 42020 71864 42076
rect 71920 42020 71944 42076
rect 72000 42020 72024 42076
rect 72080 42020 72104 42076
rect 72160 42020 72188 42076
rect 71836 41996 72188 42020
rect 71836 41940 71864 41996
rect 71920 41940 71944 41996
rect 72000 41940 72024 41996
rect 72080 41940 72104 41996
rect 72160 41940 72188 41996
rect 71836 41914 72188 41940
rect 71836 41862 71858 41914
rect 71910 41862 71922 41914
rect 71974 41862 71986 41914
rect 72038 41862 72050 41914
rect 72102 41862 72114 41914
rect 72166 41862 72188 41914
rect 71836 40826 72188 41862
rect 71836 40774 71858 40826
rect 71910 40774 71922 40826
rect 71974 40774 71986 40826
rect 72038 40774 72050 40826
rect 72102 40774 72114 40826
rect 72166 40774 72188 40826
rect 71836 39738 72188 40774
rect 71836 39686 71858 39738
rect 71910 39686 71922 39738
rect 71974 39686 71986 39738
rect 72038 39686 72050 39738
rect 72102 39686 72114 39738
rect 72166 39686 72188 39738
rect 71836 38650 72188 39686
rect 71836 38598 71858 38650
rect 71910 38598 71922 38650
rect 71974 38598 71986 38650
rect 72038 38598 72050 38650
rect 72102 38598 72114 38650
rect 72166 38598 72188 38650
rect 71836 37562 72188 38598
rect 71836 37510 71858 37562
rect 71910 37510 71922 37562
rect 71974 37510 71986 37562
rect 72038 37510 72050 37562
rect 72102 37510 72114 37562
rect 72166 37510 72188 37562
rect 71836 36474 72188 37510
rect 71836 36422 71858 36474
rect 71910 36422 71922 36474
rect 71974 36422 71986 36474
rect 72038 36422 72050 36474
rect 72102 36422 72114 36474
rect 72166 36422 72188 36474
rect 71836 35386 72188 36422
rect 71836 35334 71858 35386
rect 71910 35334 71922 35386
rect 71974 35334 71986 35386
rect 72038 35334 72050 35386
rect 72102 35334 72114 35386
rect 72166 35334 72188 35386
rect 71836 34298 72188 35334
rect 71836 34246 71858 34298
rect 71910 34246 71922 34298
rect 71974 34246 71986 34298
rect 72038 34246 72050 34298
rect 72102 34246 72114 34298
rect 72166 34246 72188 34298
rect 71836 33210 72188 34246
rect 71836 33158 71858 33210
rect 71910 33158 71922 33210
rect 71974 33158 71986 33210
rect 72038 33158 72050 33210
rect 72102 33158 72114 33210
rect 72166 33158 72188 33210
rect 71836 32236 72188 33158
rect 71836 32180 71864 32236
rect 71920 32180 71944 32236
rect 72000 32180 72024 32236
rect 72080 32180 72104 32236
rect 72160 32180 72188 32236
rect 71836 32156 72188 32180
rect 71836 32122 71864 32156
rect 71920 32122 71944 32156
rect 72000 32122 72024 32156
rect 72080 32122 72104 32156
rect 72160 32122 72188 32156
rect 71836 32070 71858 32122
rect 71920 32100 71922 32122
rect 72102 32100 72104 32122
rect 71910 32076 71922 32100
rect 71974 32076 71986 32100
rect 72038 32076 72050 32100
rect 72102 32076 72114 32100
rect 71920 32070 71922 32076
rect 72102 32070 72104 32076
rect 72166 32070 72188 32122
rect 71836 32020 71864 32070
rect 71920 32020 71944 32070
rect 72000 32020 72024 32070
rect 72080 32020 72104 32070
rect 72160 32020 72188 32070
rect 71836 31996 72188 32020
rect 71836 31940 71864 31996
rect 71920 31940 71944 31996
rect 72000 31940 72024 31996
rect 72080 31940 72104 31996
rect 72160 31940 72188 31996
rect 71836 31034 72188 31940
rect 71836 30982 71858 31034
rect 71910 30982 71922 31034
rect 71974 30982 71986 31034
rect 72038 30982 72050 31034
rect 72102 30982 72114 31034
rect 72166 30982 72188 31034
rect 71836 29946 72188 30982
rect 71836 29894 71858 29946
rect 71910 29894 71922 29946
rect 71974 29894 71986 29946
rect 72038 29894 72050 29946
rect 72102 29894 72114 29946
rect 72166 29894 72188 29946
rect 71836 28858 72188 29894
rect 71836 28806 71858 28858
rect 71910 28806 71922 28858
rect 71974 28806 71986 28858
rect 72038 28806 72050 28858
rect 72102 28806 72114 28858
rect 72166 28806 72188 28858
rect 71836 27770 72188 28806
rect 71836 27718 71858 27770
rect 71910 27718 71922 27770
rect 71974 27718 71986 27770
rect 72038 27718 72050 27770
rect 72102 27718 72114 27770
rect 72166 27718 72188 27770
rect 71836 26682 72188 27718
rect 71836 26630 71858 26682
rect 71910 26630 71922 26682
rect 71974 26630 71986 26682
rect 72038 26630 72050 26682
rect 72102 26630 72114 26682
rect 72166 26630 72188 26682
rect 71836 25594 72188 26630
rect 71836 25542 71858 25594
rect 71910 25542 71922 25594
rect 71974 25542 71986 25594
rect 72038 25542 72050 25594
rect 72102 25542 72114 25594
rect 72166 25542 72188 25594
rect 71836 24506 72188 25542
rect 71836 24454 71858 24506
rect 71910 24454 71922 24506
rect 71974 24454 71986 24506
rect 72038 24454 72050 24506
rect 72102 24454 72114 24506
rect 72166 24454 72188 24506
rect 71836 23418 72188 24454
rect 71836 23366 71858 23418
rect 71910 23366 71922 23418
rect 71974 23366 71986 23418
rect 72038 23366 72050 23418
rect 72102 23366 72114 23418
rect 72166 23366 72188 23418
rect 71836 22330 72188 23366
rect 71836 22278 71858 22330
rect 71910 22278 71922 22330
rect 71974 22278 71986 22330
rect 72038 22278 72050 22330
rect 72102 22278 72114 22330
rect 72166 22278 72188 22330
rect 71836 22236 72188 22278
rect 71836 22180 71864 22236
rect 71920 22180 71944 22236
rect 72000 22180 72024 22236
rect 72080 22180 72104 22236
rect 72160 22180 72188 22236
rect 71836 22156 72188 22180
rect 71836 22100 71864 22156
rect 71920 22100 71944 22156
rect 72000 22100 72024 22156
rect 72080 22100 72104 22156
rect 72160 22100 72188 22156
rect 71836 22076 72188 22100
rect 71836 22020 71864 22076
rect 71920 22020 71944 22076
rect 72000 22020 72024 22076
rect 72080 22020 72104 22076
rect 72160 22020 72188 22076
rect 71836 21996 72188 22020
rect 71836 21940 71864 21996
rect 71920 21940 71944 21996
rect 72000 21940 72024 21996
rect 72080 21940 72104 21996
rect 72160 21940 72188 21996
rect 71836 21242 72188 21940
rect 71836 21190 71858 21242
rect 71910 21190 71922 21242
rect 71974 21190 71986 21242
rect 72038 21190 72050 21242
rect 72102 21190 72114 21242
rect 72166 21190 72188 21242
rect 71836 20154 72188 21190
rect 71836 20102 71858 20154
rect 71910 20102 71922 20154
rect 71974 20102 71986 20154
rect 72038 20102 72050 20154
rect 72102 20102 72114 20154
rect 72166 20102 72188 20154
rect 71836 19066 72188 20102
rect 72332 19236 72384 19242
rect 72332 19178 72384 19184
rect 71836 19014 71858 19066
rect 71910 19014 71922 19066
rect 71974 19014 71986 19066
rect 72038 19014 72050 19066
rect 72102 19014 72114 19066
rect 72166 19014 72188 19066
rect 71836 17978 72188 19014
rect 71836 17926 71858 17978
rect 71910 17926 71922 17978
rect 71974 17926 71986 17978
rect 72038 17926 72050 17978
rect 72102 17926 72114 17978
rect 72166 17926 72188 17978
rect 71836 16890 72188 17926
rect 72240 17128 72292 17134
rect 72240 17070 72292 17076
rect 71836 16838 71858 16890
rect 71910 16838 71922 16890
rect 71974 16838 71986 16890
rect 72038 16838 72050 16890
rect 72102 16838 72114 16890
rect 72166 16838 72188 16890
rect 71836 15802 72188 16838
rect 71836 15750 71858 15802
rect 71910 15750 71922 15802
rect 71974 15750 71986 15802
rect 72038 15750 72050 15802
rect 72102 15750 72114 15802
rect 72166 15750 72188 15802
rect 71836 14714 72188 15750
rect 71836 14662 71858 14714
rect 71910 14662 71922 14714
rect 71974 14662 71986 14714
rect 72038 14662 72050 14714
rect 72102 14662 72114 14714
rect 72166 14662 72188 14714
rect 71836 13626 72188 14662
rect 71836 13574 71858 13626
rect 71910 13574 71922 13626
rect 71974 13574 71986 13626
rect 72038 13574 72050 13626
rect 72102 13574 72114 13626
rect 72166 13574 72188 13626
rect 71836 12538 72188 13574
rect 71836 12486 71858 12538
rect 71910 12486 71922 12538
rect 71974 12486 71986 12538
rect 72038 12486 72050 12538
rect 72102 12486 72114 12538
rect 72166 12486 72188 12538
rect 71836 12236 72188 12486
rect 71836 12180 71864 12236
rect 71920 12180 71944 12236
rect 72000 12180 72024 12236
rect 72080 12180 72104 12236
rect 72160 12180 72188 12236
rect 71836 12156 72188 12180
rect 71836 12100 71864 12156
rect 71920 12100 71944 12156
rect 72000 12100 72024 12156
rect 72080 12100 72104 12156
rect 72160 12100 72188 12156
rect 71836 12076 72188 12100
rect 71836 12020 71864 12076
rect 71920 12020 71944 12076
rect 72000 12020 72024 12076
rect 72080 12020 72104 12076
rect 72160 12020 72188 12076
rect 71836 11996 72188 12020
rect 71836 11940 71864 11996
rect 71920 11940 71944 11996
rect 72000 11940 72024 11996
rect 72080 11940 72104 11996
rect 72160 11940 72188 11996
rect 71836 11450 72188 11940
rect 71836 11398 71858 11450
rect 71910 11398 71922 11450
rect 71974 11398 71986 11450
rect 72038 11398 72050 11450
rect 72102 11398 72114 11450
rect 72166 11398 72188 11450
rect 71836 10362 72188 11398
rect 71836 10310 71858 10362
rect 71910 10310 71922 10362
rect 71974 10310 71986 10362
rect 72038 10310 72050 10362
rect 72102 10310 72114 10362
rect 72166 10310 72188 10362
rect 71836 9274 72188 10310
rect 71836 9222 71858 9274
rect 71910 9222 71922 9274
rect 71974 9222 71986 9274
rect 72038 9222 72050 9274
rect 72102 9222 72114 9274
rect 72166 9222 72188 9274
rect 71836 8186 72188 9222
rect 71836 8134 71858 8186
rect 71910 8134 71922 8186
rect 71974 8134 71986 8186
rect 72038 8134 72050 8186
rect 72102 8134 72114 8186
rect 72166 8134 72188 8186
rect 71836 7098 72188 8134
rect 71836 7046 71858 7098
rect 71910 7046 71922 7098
rect 71974 7046 71986 7098
rect 72038 7046 72050 7098
rect 72102 7046 72114 7098
rect 72166 7046 72188 7098
rect 71836 6010 72188 7046
rect 71836 5958 71858 6010
rect 71910 5958 71922 6010
rect 71974 5958 71986 6010
rect 72038 5958 72050 6010
rect 72102 5958 72114 6010
rect 72166 5958 72188 6010
rect 71836 4922 72188 5958
rect 72252 5914 72280 17070
rect 72240 5908 72292 5914
rect 72240 5850 72292 5856
rect 71836 4870 71858 4922
rect 71910 4870 71922 4922
rect 71974 4870 71986 4922
rect 72038 4870 72050 4922
rect 72102 4870 72114 4922
rect 72166 4870 72188 4922
rect 71836 3834 72188 4870
rect 71836 3782 71858 3834
rect 71910 3782 71922 3834
rect 71974 3782 71986 3834
rect 72038 3782 72050 3834
rect 72102 3782 72114 3834
rect 72166 3782 72188 3834
rect 71836 2746 72188 3782
rect 72240 2848 72292 2854
rect 72240 2790 72292 2796
rect 71836 2694 71858 2746
rect 71910 2694 71922 2746
rect 71974 2694 71986 2746
rect 72038 2694 72050 2746
rect 72102 2694 72114 2746
rect 72166 2694 72188 2746
rect 71836 2236 72188 2694
rect 72252 2514 72280 2790
rect 72240 2508 72292 2514
rect 72240 2450 72292 2456
rect 72240 2372 72292 2378
rect 72240 2314 72292 2320
rect 71836 2180 71864 2236
rect 71920 2180 71944 2236
rect 72000 2180 72024 2236
rect 72080 2180 72104 2236
rect 72160 2180 72188 2236
rect 71836 2156 72188 2180
rect 71836 2100 71864 2156
rect 71920 2100 71944 2156
rect 72000 2100 72024 2156
rect 72080 2100 72104 2156
rect 72160 2100 72188 2156
rect 71836 2076 72188 2100
rect 71836 2020 71864 2076
rect 71920 2020 71944 2076
rect 72000 2020 72024 2076
rect 72080 2020 72104 2076
rect 72160 2020 72188 2076
rect 71836 1996 72188 2020
rect 71688 1964 71740 1970
rect 71688 1906 71740 1912
rect 71836 1940 71864 1996
rect 71920 1940 71944 1996
rect 72000 1940 72024 1996
rect 72080 1940 72104 1996
rect 72160 1940 72188 1996
rect 71320 1896 71372 1902
rect 71320 1838 71372 1844
rect 70952 1828 71004 1834
rect 70952 1770 71004 1776
rect 70768 1352 70820 1358
rect 70768 1294 70820 1300
rect 70860 1284 70912 1290
rect 70860 1226 70912 1232
rect 70872 800 70900 1226
rect 71332 800 71360 1838
rect 71836 1658 72188 1940
rect 71836 1606 71858 1658
rect 71910 1606 71922 1658
rect 71974 1606 71986 1658
rect 72038 1606 72050 1658
rect 72102 1606 72114 1658
rect 72166 1606 72188 1658
rect 71836 1040 72188 1606
rect 72252 1358 72280 2314
rect 72344 2106 72372 19178
rect 72424 18760 72476 18766
rect 72424 18702 72476 18708
rect 72436 3534 72464 18702
rect 72516 16652 72568 16658
rect 72516 16594 72568 16600
rect 72424 3528 72476 3534
rect 72424 3470 72476 3476
rect 72528 3398 72556 16594
rect 72608 14884 72660 14890
rect 72608 14826 72660 14832
rect 72516 3392 72568 3398
rect 72516 3334 72568 3340
rect 72332 2100 72384 2106
rect 72332 2042 72384 2048
rect 72240 1352 72292 1358
rect 72240 1294 72292 1300
rect 72620 950 72648 14826
rect 72700 3052 72752 3058
rect 72700 2994 72752 3000
rect 72712 1358 72740 2994
rect 72700 1352 72752 1358
rect 72700 1294 72752 1300
rect 72608 944 72660 950
rect 72608 886 72660 892
rect 70492 740 70544 746
rect 70492 682 70544 688
rect 70858 0 70914 800
rect 71318 0 71374 800
rect 72804 406 72832 67730
rect 74188 67482 74540 68518
rect 74188 67430 74210 67482
rect 74262 67430 74274 67482
rect 74326 67430 74338 67482
rect 74390 67430 74402 67482
rect 74454 67430 74466 67482
rect 74518 67430 74540 67482
rect 74188 66394 74540 67430
rect 74188 66342 74210 66394
rect 74262 66342 74274 66394
rect 74326 66342 74338 66394
rect 74390 66342 74402 66394
rect 74454 66342 74466 66394
rect 74518 66342 74540 66394
rect 74188 65306 74540 66342
rect 74188 65254 74210 65306
rect 74262 65254 74274 65306
rect 74326 65254 74338 65306
rect 74390 65254 74402 65306
rect 74454 65254 74466 65306
rect 74518 65254 74540 65306
rect 74188 64588 74540 65254
rect 74188 64532 74216 64588
rect 74272 64532 74296 64588
rect 74352 64532 74376 64588
rect 74432 64532 74456 64588
rect 74512 64532 74540 64588
rect 74188 64508 74540 64532
rect 74188 64452 74216 64508
rect 74272 64452 74296 64508
rect 74352 64452 74376 64508
rect 74432 64452 74456 64508
rect 74512 64452 74540 64508
rect 74188 64428 74540 64452
rect 74188 64372 74216 64428
rect 74272 64372 74296 64428
rect 74352 64372 74376 64428
rect 74432 64372 74456 64428
rect 74512 64372 74540 64428
rect 74188 64348 74540 64372
rect 74188 64292 74216 64348
rect 74272 64292 74296 64348
rect 74352 64292 74376 64348
rect 74432 64292 74456 64348
rect 74512 64292 74540 64348
rect 74188 64218 74540 64292
rect 74188 64166 74210 64218
rect 74262 64166 74274 64218
rect 74326 64166 74338 64218
rect 74390 64166 74402 64218
rect 74454 64166 74466 64218
rect 74518 64166 74540 64218
rect 74188 63130 74540 64166
rect 74188 63078 74210 63130
rect 74262 63078 74274 63130
rect 74326 63078 74338 63130
rect 74390 63078 74402 63130
rect 74454 63078 74466 63130
rect 74518 63078 74540 63130
rect 74188 62042 74540 63078
rect 74188 61990 74210 62042
rect 74262 61990 74274 62042
rect 74326 61990 74338 62042
rect 74390 61990 74402 62042
rect 74454 61990 74466 62042
rect 74518 61990 74540 62042
rect 74188 60954 74540 61990
rect 74188 60902 74210 60954
rect 74262 60902 74274 60954
rect 74326 60902 74338 60954
rect 74390 60902 74402 60954
rect 74454 60902 74466 60954
rect 74518 60902 74540 60954
rect 74188 59866 74540 60902
rect 74188 59814 74210 59866
rect 74262 59814 74274 59866
rect 74326 59814 74338 59866
rect 74390 59814 74402 59866
rect 74454 59814 74466 59866
rect 74518 59814 74540 59866
rect 74188 58778 74540 59814
rect 74188 58726 74210 58778
rect 74262 58726 74274 58778
rect 74326 58726 74338 58778
rect 74390 58726 74402 58778
rect 74454 58726 74466 58778
rect 74518 58726 74540 58778
rect 74188 57690 74540 58726
rect 74188 57638 74210 57690
rect 74262 57638 74274 57690
rect 74326 57638 74338 57690
rect 74390 57638 74402 57690
rect 74454 57638 74466 57690
rect 74518 57638 74540 57690
rect 74188 56602 74540 57638
rect 74188 56550 74210 56602
rect 74262 56550 74274 56602
rect 74326 56550 74338 56602
rect 74390 56550 74402 56602
rect 74454 56550 74466 56602
rect 74518 56550 74540 56602
rect 74188 55514 74540 56550
rect 74188 55462 74210 55514
rect 74262 55462 74274 55514
rect 74326 55462 74338 55514
rect 74390 55462 74402 55514
rect 74454 55462 74466 55514
rect 74518 55462 74540 55514
rect 74188 54588 74540 55462
rect 74188 54532 74216 54588
rect 74272 54532 74296 54588
rect 74352 54532 74376 54588
rect 74432 54532 74456 54588
rect 74512 54532 74540 54588
rect 74188 54508 74540 54532
rect 74188 54452 74216 54508
rect 74272 54452 74296 54508
rect 74352 54452 74376 54508
rect 74432 54452 74456 54508
rect 74512 54452 74540 54508
rect 74188 54428 74540 54452
rect 74188 54426 74216 54428
rect 74272 54426 74296 54428
rect 74352 54426 74376 54428
rect 74432 54426 74456 54428
rect 74512 54426 74540 54428
rect 74188 54374 74210 54426
rect 74272 54374 74274 54426
rect 74454 54374 74456 54426
rect 74518 54374 74540 54426
rect 74188 54372 74216 54374
rect 74272 54372 74296 54374
rect 74352 54372 74376 54374
rect 74432 54372 74456 54374
rect 74512 54372 74540 54374
rect 74188 54348 74540 54372
rect 74188 54292 74216 54348
rect 74272 54292 74296 54348
rect 74352 54292 74376 54348
rect 74432 54292 74456 54348
rect 74512 54292 74540 54348
rect 74188 53338 74540 54292
rect 74188 53286 74210 53338
rect 74262 53286 74274 53338
rect 74326 53286 74338 53338
rect 74390 53286 74402 53338
rect 74454 53286 74466 53338
rect 74518 53286 74540 53338
rect 74188 52250 74540 53286
rect 74188 52198 74210 52250
rect 74262 52198 74274 52250
rect 74326 52198 74338 52250
rect 74390 52198 74402 52250
rect 74454 52198 74466 52250
rect 74518 52198 74540 52250
rect 74188 51162 74540 52198
rect 74188 51110 74210 51162
rect 74262 51110 74274 51162
rect 74326 51110 74338 51162
rect 74390 51110 74402 51162
rect 74454 51110 74466 51162
rect 74518 51110 74540 51162
rect 74188 50074 74540 51110
rect 74188 50022 74210 50074
rect 74262 50022 74274 50074
rect 74326 50022 74338 50074
rect 74390 50022 74402 50074
rect 74454 50022 74466 50074
rect 74518 50022 74540 50074
rect 74188 48986 74540 50022
rect 74188 48934 74210 48986
rect 74262 48934 74274 48986
rect 74326 48934 74338 48986
rect 74390 48934 74402 48986
rect 74454 48934 74466 48986
rect 74518 48934 74540 48986
rect 74188 47898 74540 48934
rect 74188 47846 74210 47898
rect 74262 47846 74274 47898
rect 74326 47846 74338 47898
rect 74390 47846 74402 47898
rect 74454 47846 74466 47898
rect 74518 47846 74540 47898
rect 74188 46810 74540 47846
rect 74188 46758 74210 46810
rect 74262 46758 74274 46810
rect 74326 46758 74338 46810
rect 74390 46758 74402 46810
rect 74454 46758 74466 46810
rect 74518 46758 74540 46810
rect 74188 45722 74540 46758
rect 74188 45670 74210 45722
rect 74262 45670 74274 45722
rect 74326 45670 74338 45722
rect 74390 45670 74402 45722
rect 74454 45670 74466 45722
rect 74518 45670 74540 45722
rect 74188 44634 74540 45670
rect 74188 44582 74210 44634
rect 74262 44588 74274 44634
rect 74326 44588 74338 44634
rect 74390 44588 74402 44634
rect 74454 44588 74466 44634
rect 74272 44582 74274 44588
rect 74454 44582 74456 44588
rect 74518 44582 74540 44634
rect 74188 44532 74216 44582
rect 74272 44532 74296 44582
rect 74352 44532 74376 44582
rect 74432 44532 74456 44582
rect 74512 44532 74540 44582
rect 74188 44508 74540 44532
rect 74188 44452 74216 44508
rect 74272 44452 74296 44508
rect 74352 44452 74376 44508
rect 74432 44452 74456 44508
rect 74512 44452 74540 44508
rect 74188 44428 74540 44452
rect 74188 44372 74216 44428
rect 74272 44372 74296 44428
rect 74352 44372 74376 44428
rect 74432 44372 74456 44428
rect 74512 44372 74540 44428
rect 74188 44348 74540 44372
rect 74188 44292 74216 44348
rect 74272 44292 74296 44348
rect 74352 44292 74376 44348
rect 74432 44292 74456 44348
rect 74512 44292 74540 44348
rect 74188 43546 74540 44292
rect 74188 43494 74210 43546
rect 74262 43494 74274 43546
rect 74326 43494 74338 43546
rect 74390 43494 74402 43546
rect 74454 43494 74466 43546
rect 74518 43494 74540 43546
rect 74188 42458 74540 43494
rect 74188 42406 74210 42458
rect 74262 42406 74274 42458
rect 74326 42406 74338 42458
rect 74390 42406 74402 42458
rect 74454 42406 74466 42458
rect 74518 42406 74540 42458
rect 74188 41370 74540 42406
rect 74188 41318 74210 41370
rect 74262 41318 74274 41370
rect 74326 41318 74338 41370
rect 74390 41318 74402 41370
rect 74454 41318 74466 41370
rect 74518 41318 74540 41370
rect 74188 40282 74540 41318
rect 74188 40230 74210 40282
rect 74262 40230 74274 40282
rect 74326 40230 74338 40282
rect 74390 40230 74402 40282
rect 74454 40230 74466 40282
rect 74518 40230 74540 40282
rect 74188 39194 74540 40230
rect 74188 39142 74210 39194
rect 74262 39142 74274 39194
rect 74326 39142 74338 39194
rect 74390 39142 74402 39194
rect 74454 39142 74466 39194
rect 74518 39142 74540 39194
rect 74188 38106 74540 39142
rect 74188 38054 74210 38106
rect 74262 38054 74274 38106
rect 74326 38054 74338 38106
rect 74390 38054 74402 38106
rect 74454 38054 74466 38106
rect 74518 38054 74540 38106
rect 74188 37018 74540 38054
rect 74188 36966 74210 37018
rect 74262 36966 74274 37018
rect 74326 36966 74338 37018
rect 74390 36966 74402 37018
rect 74454 36966 74466 37018
rect 74518 36966 74540 37018
rect 74188 35930 74540 36966
rect 74188 35878 74210 35930
rect 74262 35878 74274 35930
rect 74326 35878 74338 35930
rect 74390 35878 74402 35930
rect 74454 35878 74466 35930
rect 74518 35878 74540 35930
rect 74188 34842 74540 35878
rect 74188 34790 74210 34842
rect 74262 34790 74274 34842
rect 74326 34790 74338 34842
rect 74390 34790 74402 34842
rect 74454 34790 74466 34842
rect 74518 34790 74540 34842
rect 74188 34588 74540 34790
rect 74188 34532 74216 34588
rect 74272 34532 74296 34588
rect 74352 34532 74376 34588
rect 74432 34532 74456 34588
rect 74512 34532 74540 34588
rect 74188 34508 74540 34532
rect 74188 34452 74216 34508
rect 74272 34452 74296 34508
rect 74352 34452 74376 34508
rect 74432 34452 74456 34508
rect 74512 34452 74540 34508
rect 74188 34428 74540 34452
rect 74188 34372 74216 34428
rect 74272 34372 74296 34428
rect 74352 34372 74376 34428
rect 74432 34372 74456 34428
rect 74512 34372 74540 34428
rect 74188 34348 74540 34372
rect 74188 34292 74216 34348
rect 74272 34292 74296 34348
rect 74352 34292 74376 34348
rect 74432 34292 74456 34348
rect 74512 34292 74540 34348
rect 74188 33754 74540 34292
rect 74188 33702 74210 33754
rect 74262 33702 74274 33754
rect 74326 33702 74338 33754
rect 74390 33702 74402 33754
rect 74454 33702 74466 33754
rect 74518 33702 74540 33754
rect 74188 32666 74540 33702
rect 74188 32614 74210 32666
rect 74262 32614 74274 32666
rect 74326 32614 74338 32666
rect 74390 32614 74402 32666
rect 74454 32614 74466 32666
rect 74518 32614 74540 32666
rect 74188 31578 74540 32614
rect 74188 31526 74210 31578
rect 74262 31526 74274 31578
rect 74326 31526 74338 31578
rect 74390 31526 74402 31578
rect 74454 31526 74466 31578
rect 74518 31526 74540 31578
rect 74188 30490 74540 31526
rect 74188 30438 74210 30490
rect 74262 30438 74274 30490
rect 74326 30438 74338 30490
rect 74390 30438 74402 30490
rect 74454 30438 74466 30490
rect 74518 30438 74540 30490
rect 74188 29402 74540 30438
rect 74188 29350 74210 29402
rect 74262 29350 74274 29402
rect 74326 29350 74338 29402
rect 74390 29350 74402 29402
rect 74454 29350 74466 29402
rect 74518 29350 74540 29402
rect 74188 28314 74540 29350
rect 74188 28262 74210 28314
rect 74262 28262 74274 28314
rect 74326 28262 74338 28314
rect 74390 28262 74402 28314
rect 74454 28262 74466 28314
rect 74518 28262 74540 28314
rect 74188 27226 74540 28262
rect 74188 27174 74210 27226
rect 74262 27174 74274 27226
rect 74326 27174 74338 27226
rect 74390 27174 74402 27226
rect 74454 27174 74466 27226
rect 74518 27174 74540 27226
rect 74188 26138 74540 27174
rect 74188 26086 74210 26138
rect 74262 26086 74274 26138
rect 74326 26086 74338 26138
rect 74390 26086 74402 26138
rect 74454 26086 74466 26138
rect 74518 26086 74540 26138
rect 74188 25050 74540 26086
rect 74188 24998 74210 25050
rect 74262 24998 74274 25050
rect 74326 24998 74338 25050
rect 74390 24998 74402 25050
rect 74454 24998 74466 25050
rect 74518 24998 74540 25050
rect 74188 24588 74540 24998
rect 74188 24532 74216 24588
rect 74272 24532 74296 24588
rect 74352 24532 74376 24588
rect 74432 24532 74456 24588
rect 74512 24532 74540 24588
rect 74188 24508 74540 24532
rect 74188 24452 74216 24508
rect 74272 24452 74296 24508
rect 74352 24452 74376 24508
rect 74432 24452 74456 24508
rect 74512 24452 74540 24508
rect 74188 24428 74540 24452
rect 74188 24372 74216 24428
rect 74272 24372 74296 24428
rect 74352 24372 74376 24428
rect 74432 24372 74456 24428
rect 74512 24372 74540 24428
rect 74188 24348 74540 24372
rect 74188 24292 74216 24348
rect 74272 24292 74296 24348
rect 74352 24292 74376 24348
rect 74432 24292 74456 24348
rect 74512 24292 74540 24348
rect 74188 23962 74540 24292
rect 74188 23910 74210 23962
rect 74262 23910 74274 23962
rect 74326 23910 74338 23962
rect 74390 23910 74402 23962
rect 74454 23910 74466 23962
rect 74518 23910 74540 23962
rect 74188 22874 74540 23910
rect 74188 22822 74210 22874
rect 74262 22822 74274 22874
rect 74326 22822 74338 22874
rect 74390 22822 74402 22874
rect 74454 22822 74466 22874
rect 74518 22822 74540 22874
rect 74188 21786 74540 22822
rect 74188 21734 74210 21786
rect 74262 21734 74274 21786
rect 74326 21734 74338 21786
rect 74390 21734 74402 21786
rect 74454 21734 74466 21786
rect 74518 21734 74540 21786
rect 74188 20698 74540 21734
rect 74188 20646 74210 20698
rect 74262 20646 74274 20698
rect 74326 20646 74338 20698
rect 74390 20646 74402 20698
rect 74454 20646 74466 20698
rect 74518 20646 74540 20698
rect 74188 19610 74540 20646
rect 74188 19558 74210 19610
rect 74262 19558 74274 19610
rect 74326 19558 74338 19610
rect 74390 19558 74402 19610
rect 74454 19558 74466 19610
rect 74518 19558 74540 19610
rect 74188 18522 74540 19558
rect 74188 18470 74210 18522
rect 74262 18470 74274 18522
rect 74326 18470 74338 18522
rect 74390 18470 74402 18522
rect 74454 18470 74466 18522
rect 74518 18470 74540 18522
rect 74188 17434 74540 18470
rect 74188 17382 74210 17434
rect 74262 17382 74274 17434
rect 74326 17382 74338 17434
rect 74390 17382 74402 17434
rect 74454 17382 74466 17434
rect 74518 17382 74540 17434
rect 74188 16346 74540 17382
rect 74188 16294 74210 16346
rect 74262 16294 74274 16346
rect 74326 16294 74338 16346
rect 74390 16294 74402 16346
rect 74454 16294 74466 16346
rect 74518 16294 74540 16346
rect 74188 15258 74540 16294
rect 74188 15206 74210 15258
rect 74262 15206 74274 15258
rect 74326 15206 74338 15258
rect 74390 15206 74402 15258
rect 74454 15206 74466 15258
rect 74518 15206 74540 15258
rect 74188 14588 74540 15206
rect 74188 14532 74216 14588
rect 74272 14532 74296 14588
rect 74352 14532 74376 14588
rect 74432 14532 74456 14588
rect 74512 14532 74540 14588
rect 74188 14508 74540 14532
rect 74188 14452 74216 14508
rect 74272 14452 74296 14508
rect 74352 14452 74376 14508
rect 74432 14452 74456 14508
rect 74512 14452 74540 14508
rect 74188 14428 74540 14452
rect 74188 14372 74216 14428
rect 74272 14372 74296 14428
rect 74352 14372 74376 14428
rect 74432 14372 74456 14428
rect 74512 14372 74540 14428
rect 74188 14348 74540 14372
rect 74188 14292 74216 14348
rect 74272 14292 74296 14348
rect 74352 14292 74376 14348
rect 74432 14292 74456 14348
rect 74512 14292 74540 14348
rect 74188 14170 74540 14292
rect 74188 14118 74210 14170
rect 74262 14118 74274 14170
rect 74326 14118 74338 14170
rect 74390 14118 74402 14170
rect 74454 14118 74466 14170
rect 74518 14118 74540 14170
rect 74188 13082 74540 14118
rect 74188 13030 74210 13082
rect 74262 13030 74274 13082
rect 74326 13030 74338 13082
rect 74390 13030 74402 13082
rect 74454 13030 74466 13082
rect 74518 13030 74540 13082
rect 74188 11994 74540 13030
rect 74188 11942 74210 11994
rect 74262 11942 74274 11994
rect 74326 11942 74338 11994
rect 74390 11942 74402 11994
rect 74454 11942 74466 11994
rect 74518 11942 74540 11994
rect 74188 10906 74540 11942
rect 74188 10854 74210 10906
rect 74262 10854 74274 10906
rect 74326 10854 74338 10906
rect 74390 10854 74402 10906
rect 74454 10854 74466 10906
rect 74518 10854 74540 10906
rect 74188 9818 74540 10854
rect 74188 9766 74210 9818
rect 74262 9766 74274 9818
rect 74326 9766 74338 9818
rect 74390 9766 74402 9818
rect 74454 9766 74466 9818
rect 74518 9766 74540 9818
rect 74188 8730 74540 9766
rect 74188 8678 74210 8730
rect 74262 8678 74274 8730
rect 74326 8678 74338 8730
rect 74390 8678 74402 8730
rect 74454 8678 74466 8730
rect 74518 8678 74540 8730
rect 74188 7642 74540 8678
rect 74188 7590 74210 7642
rect 74262 7590 74274 7642
rect 74326 7590 74338 7642
rect 74390 7590 74402 7642
rect 74454 7590 74466 7642
rect 74518 7590 74540 7642
rect 74188 6554 74540 7590
rect 74188 6502 74210 6554
rect 74262 6502 74274 6554
rect 74326 6502 74338 6554
rect 74390 6502 74402 6554
rect 74454 6502 74466 6554
rect 74518 6502 74540 6554
rect 73436 5568 73488 5574
rect 73436 5510 73488 5516
rect 73252 2984 73304 2990
rect 73252 2926 73304 2932
rect 73264 1358 73292 2926
rect 73448 2038 73476 5510
rect 74188 5466 74540 6502
rect 74188 5414 74210 5466
rect 74262 5414 74274 5466
rect 74326 5414 74338 5466
rect 74390 5414 74402 5466
rect 74454 5414 74466 5466
rect 74518 5414 74540 5466
rect 74188 4588 74540 5414
rect 74188 4532 74216 4588
rect 74272 4532 74296 4588
rect 74352 4532 74376 4588
rect 74432 4532 74456 4588
rect 74512 4532 74540 4588
rect 74188 4508 74540 4532
rect 74188 4452 74216 4508
rect 74272 4452 74296 4508
rect 74352 4452 74376 4508
rect 74432 4452 74456 4508
rect 74512 4452 74540 4508
rect 74188 4428 74540 4452
rect 74188 4378 74216 4428
rect 74272 4378 74296 4428
rect 74352 4378 74376 4428
rect 74432 4378 74456 4428
rect 74512 4378 74540 4428
rect 74188 4326 74210 4378
rect 74272 4372 74274 4378
rect 74454 4372 74456 4378
rect 74262 4348 74274 4372
rect 74326 4348 74338 4372
rect 74390 4348 74402 4372
rect 74454 4348 74466 4372
rect 74272 4326 74274 4348
rect 74454 4326 74456 4348
rect 74518 4326 74540 4378
rect 74188 4292 74216 4326
rect 74272 4292 74296 4326
rect 74352 4292 74376 4326
rect 74432 4292 74456 4326
rect 74512 4292 74540 4326
rect 74188 3290 74540 4292
rect 74188 3238 74210 3290
rect 74262 3238 74274 3290
rect 74326 3238 74338 3290
rect 74390 3238 74402 3290
rect 74454 3238 74466 3290
rect 74518 3238 74540 3290
rect 74188 2202 74540 3238
rect 74632 2304 74684 2310
rect 74632 2246 74684 2252
rect 74188 2150 74210 2202
rect 74262 2150 74274 2202
rect 74326 2150 74338 2202
rect 74390 2150 74402 2202
rect 74454 2150 74466 2202
rect 74518 2150 74540 2202
rect 73436 2032 73488 2038
rect 73436 1974 73488 1980
rect 73712 1964 73764 1970
rect 73712 1906 73764 1912
rect 73724 1562 73752 1906
rect 73712 1556 73764 1562
rect 73712 1498 73764 1504
rect 73252 1352 73304 1358
rect 73252 1294 73304 1300
rect 74188 1114 74540 2150
rect 74644 1426 74672 2246
rect 74632 1420 74684 1426
rect 74632 1362 74684 1368
rect 74188 1062 74210 1114
rect 74262 1062 74274 1114
rect 74326 1062 74338 1114
rect 74390 1062 74402 1114
rect 74454 1062 74466 1114
rect 74518 1062 74540 1114
rect 74188 1040 74540 1062
rect 72792 400 72844 406
rect 72792 342 72844 348
<< via2 >>
rect 2044 84532 2100 84588
rect 2044 84452 2100 84508
rect 2044 84372 2100 84428
rect 2044 84292 2100 84348
rect 5540 84532 5596 84588
rect 5540 84452 5596 84508
rect 5540 84372 5596 84428
rect 5540 84292 5596 84348
rect 8430 84532 8486 84588
rect 8430 84452 8486 84508
rect 8430 84372 8486 84428
rect 8430 84292 8486 84348
rect 11320 84532 11376 84588
rect 11320 84452 11376 84508
rect 11320 84372 11376 84428
rect 11320 84292 11376 84348
rect 14210 84532 14266 84588
rect 14210 84452 14266 84508
rect 14210 84372 14266 84428
rect 14210 84292 14266 84348
rect 17100 84532 17156 84588
rect 17100 84452 17156 84508
rect 17100 84372 17156 84428
rect 17100 84292 17156 84348
rect 19990 84532 20046 84588
rect 19990 84452 20046 84508
rect 19990 84372 20046 84428
rect 19990 84292 20046 84348
rect 22880 84532 22936 84588
rect 22880 84452 22936 84508
rect 22880 84372 22936 84428
rect 22880 84292 22936 84348
rect 25770 84532 25826 84588
rect 25770 84452 25826 84508
rect 25770 84372 25826 84428
rect 25770 84292 25826 84348
rect 28660 84532 28716 84588
rect 28660 84452 28716 84508
rect 28660 84372 28716 84428
rect 28660 84292 28716 84348
rect 31550 84532 31606 84588
rect 31550 84452 31606 84508
rect 31550 84372 31606 84428
rect 31550 84292 31606 84348
rect 34440 84532 34496 84588
rect 34440 84452 34496 84508
rect 34440 84372 34496 84428
rect 34440 84292 34496 84348
rect 37330 84532 37386 84588
rect 37330 84452 37386 84508
rect 37330 84372 37386 84428
rect 37330 84292 37386 84348
rect 40220 84532 40276 84588
rect 40220 84452 40276 84508
rect 40220 84372 40276 84428
rect 40220 84292 40276 84348
rect 43110 84532 43166 84588
rect 43110 84452 43166 84508
rect 43110 84372 43166 84428
rect 43110 84292 43166 84348
rect 46000 84532 46056 84588
rect 46000 84452 46056 84508
rect 46000 84372 46056 84428
rect 46000 84292 46056 84348
rect 49008 84532 49064 84588
rect 49008 84452 49064 84508
rect 49008 84372 49064 84428
rect 49008 84292 49064 84348
rect 52237 84532 52293 84588
rect 52237 84452 52293 84508
rect 52237 84372 52293 84428
rect 52237 84292 52293 84348
rect 53638 84532 53694 84588
rect 53638 84452 53694 84508
rect 53638 84372 53694 84428
rect 53638 84292 53694 84348
rect 53806 84532 53862 84588
rect 53806 84452 53862 84508
rect 53806 84372 53862 84428
rect 53806 84292 53862 84348
rect 54550 84532 54606 84588
rect 54550 84452 54606 84508
rect 54550 84372 54606 84428
rect 54550 84292 54606 84348
rect 54940 84532 54996 84588
rect 54940 84452 54996 84508
rect 54940 84372 54996 84428
rect 54940 84292 54996 84348
rect 55656 84532 55712 84588
rect 55656 84452 55712 84508
rect 55656 84372 55712 84428
rect 55656 84292 55712 84348
rect 56234 84532 56290 84588
rect 56234 84452 56290 84508
rect 56234 84372 56290 84428
rect 56234 84292 56290 84348
rect 56679 84532 56735 84588
rect 56679 84452 56735 84508
rect 56679 84372 56735 84428
rect 56679 84292 56735 84348
rect 56983 84532 57039 84588
rect 56983 84452 57039 84508
rect 56983 84372 57039 84428
rect 56983 84292 57039 84348
rect 57825 84532 57881 84588
rect 57825 84452 57881 84508
rect 57825 84372 57881 84428
rect 57825 84292 57881 84348
rect 58465 84532 58521 84588
rect 58465 84452 58521 84508
rect 58465 84372 58521 84428
rect 58465 84292 58521 84348
rect 59048 84532 59104 84588
rect 59048 84452 59104 84508
rect 59048 84372 59104 84428
rect 59048 84292 59104 84348
rect 60326 84532 60382 84588
rect 60326 84452 60382 84508
rect 60326 84372 60382 84428
rect 60326 84292 60382 84348
rect 60484 84532 60540 84588
rect 60484 84452 60540 84508
rect 60484 84372 60540 84428
rect 60484 84292 60540 84348
rect 62528 84532 62584 84588
rect 62608 84532 62664 84588
rect 62528 84452 62584 84508
rect 62608 84452 62664 84508
rect 62528 84372 62584 84428
rect 62608 84372 62664 84428
rect 62528 84292 62584 84348
rect 62608 84292 62664 84348
rect 2184 82180 2240 82236
rect 2264 82180 2320 82236
rect 2184 82100 2240 82156
rect 2264 82100 2320 82156
rect 2184 82020 2240 82076
rect 2264 82020 2320 82076
rect 2184 81940 2240 81996
rect 2264 81940 2320 81996
rect 5393 82180 5449 82236
rect 5393 82100 5449 82156
rect 5393 82020 5449 82076
rect 5393 81940 5449 81996
rect 8283 82180 8339 82236
rect 8283 82100 8339 82156
rect 8283 82020 8339 82076
rect 8283 81940 8339 81996
rect 11173 82180 11229 82236
rect 11173 82100 11229 82156
rect 11173 82020 11229 82076
rect 11173 81940 11229 81996
rect 14063 82180 14119 82236
rect 14063 82100 14119 82156
rect 14063 82020 14119 82076
rect 14063 81940 14119 81996
rect 16953 82180 17009 82236
rect 16953 82100 17009 82156
rect 16953 82020 17009 82076
rect 16953 81940 17009 81996
rect 19843 82180 19899 82236
rect 19843 82100 19899 82156
rect 19843 82020 19899 82076
rect 19843 81940 19899 81996
rect 22733 82180 22789 82236
rect 22733 82100 22789 82156
rect 22733 82020 22789 82076
rect 22733 81940 22789 81996
rect 25623 82180 25679 82236
rect 25623 82100 25679 82156
rect 25623 82020 25679 82076
rect 25623 81940 25679 81996
rect 28513 82180 28569 82236
rect 28513 82100 28569 82156
rect 28513 82020 28569 82076
rect 28513 81940 28569 81996
rect 31403 82180 31459 82236
rect 31403 82100 31459 82156
rect 31403 82020 31459 82076
rect 31403 81940 31459 81996
rect 34293 82180 34349 82236
rect 34293 82100 34349 82156
rect 34293 82020 34349 82076
rect 34293 81940 34349 81996
rect 37183 82180 37239 82236
rect 37183 82100 37239 82156
rect 37183 82020 37239 82076
rect 37183 81940 37239 81996
rect 40073 82180 40129 82236
rect 40073 82100 40129 82156
rect 40073 82020 40129 82076
rect 40073 81940 40129 81996
rect 42963 82180 43019 82236
rect 42963 82100 43019 82156
rect 42963 82020 43019 82076
rect 42963 81940 43019 81996
rect 45853 82180 45909 82236
rect 45853 82100 45909 82156
rect 45853 82020 45909 82076
rect 45853 81940 45909 81996
rect 48800 82180 48856 82236
rect 48800 82100 48856 82156
rect 48800 82020 48856 82076
rect 48800 81940 48856 81996
rect 49662 82180 49718 82236
rect 49742 82180 49798 82236
rect 49662 82100 49718 82156
rect 49742 82100 49798 82156
rect 49662 82020 49718 82076
rect 49742 82020 49798 82076
rect 49662 81940 49718 81996
rect 49742 81940 49798 81996
rect 52956 82180 53012 82236
rect 52956 82100 53012 82156
rect 52956 82020 53012 82076
rect 52956 81940 53012 81996
rect 53114 82180 53170 82236
rect 53114 82100 53170 82156
rect 53114 82020 53170 82076
rect 53114 81940 53170 81996
rect 53470 82180 53526 82236
rect 53470 82100 53526 82156
rect 53470 82020 53526 82076
rect 53470 81940 53526 81996
rect 54788 82180 54844 82236
rect 54788 82100 54844 82156
rect 54788 82020 54844 82076
rect 54788 81940 54844 81996
rect 55381 82180 55437 82236
rect 55381 82100 55437 82156
rect 55381 82020 55437 82076
rect 55381 81940 55437 81996
rect 56527 82180 56583 82236
rect 56527 82100 56583 82156
rect 56527 82020 56583 82076
rect 56527 81940 56583 81996
rect 57963 82180 58019 82236
rect 58043 82180 58099 82236
rect 57963 82100 58019 82156
rect 58043 82100 58099 82156
rect 57963 82020 58019 82076
rect 58043 82020 58099 82076
rect 57963 81940 58019 81996
rect 58043 81940 58099 81996
rect 59206 82180 59262 82236
rect 59206 82100 59262 82156
rect 59206 82020 59262 82076
rect 59206 81940 59262 81996
rect 59364 82180 59420 82236
rect 59364 82100 59420 82156
rect 59364 82020 59420 82076
rect 59364 81940 59420 81996
rect 59672 82180 59728 82236
rect 59672 82100 59728 82156
rect 59672 82020 59728 82076
rect 59672 81940 59728 81996
rect 59818 82180 59874 82236
rect 59818 82100 59874 82156
rect 59818 82020 59874 82076
rect 59818 81940 59874 81996
rect 59954 82180 60010 82236
rect 60034 82180 60090 82236
rect 59954 82100 60010 82156
rect 60034 82100 60090 82156
rect 59954 82020 60010 82076
rect 60034 82020 60090 82076
rect 59954 81940 60010 81996
rect 60034 81940 60090 81996
rect 62326 82180 62382 82236
rect 62406 82180 62462 82236
rect 62326 82100 62382 82156
rect 62406 82100 62462 82156
rect 62326 82020 62382 82076
rect 62406 82020 62462 82076
rect 62326 81940 62382 81996
rect 62406 81940 62462 81996
rect 2044 74532 2100 74588
rect 2044 74452 2100 74508
rect 2044 74372 2100 74428
rect 2044 74292 2100 74348
rect 5540 74532 5596 74588
rect 5540 74452 5596 74508
rect 5540 74372 5596 74428
rect 5540 74292 5596 74348
rect 8430 74532 8486 74588
rect 8430 74452 8486 74508
rect 8430 74372 8486 74428
rect 8430 74292 8486 74348
rect 11320 74532 11376 74588
rect 11320 74452 11376 74508
rect 11320 74372 11376 74428
rect 11320 74292 11376 74348
rect 14210 74532 14266 74588
rect 14210 74452 14266 74508
rect 14210 74372 14266 74428
rect 14210 74292 14266 74348
rect 17100 74532 17156 74588
rect 17100 74452 17156 74508
rect 17100 74372 17156 74428
rect 17100 74292 17156 74348
rect 19990 74532 20046 74588
rect 19990 74452 20046 74508
rect 19990 74372 20046 74428
rect 19990 74292 20046 74348
rect 22880 74532 22936 74588
rect 22880 74452 22936 74508
rect 22880 74372 22936 74428
rect 22880 74292 22936 74348
rect 25770 74532 25826 74588
rect 25770 74452 25826 74508
rect 25770 74372 25826 74428
rect 25770 74292 25826 74348
rect 28660 74532 28716 74588
rect 28660 74452 28716 74508
rect 28660 74372 28716 74428
rect 28660 74292 28716 74348
rect 31550 74532 31606 74588
rect 31550 74452 31606 74508
rect 31550 74372 31606 74428
rect 31550 74292 31606 74348
rect 34440 74532 34496 74588
rect 34440 74452 34496 74508
rect 34440 74372 34496 74428
rect 34440 74292 34496 74348
rect 37330 74532 37386 74588
rect 37330 74452 37386 74508
rect 37330 74372 37386 74428
rect 37330 74292 37386 74348
rect 40220 74532 40276 74588
rect 40220 74452 40276 74508
rect 40220 74372 40276 74428
rect 40220 74292 40276 74348
rect 43110 74532 43166 74588
rect 43110 74452 43166 74508
rect 43110 74372 43166 74428
rect 43110 74292 43166 74348
rect 46000 74532 46056 74588
rect 46000 74452 46056 74508
rect 46000 74372 46056 74428
rect 46000 74292 46056 74348
rect 49008 74532 49064 74588
rect 49008 74452 49064 74508
rect 49008 74372 49064 74428
rect 49008 74292 49064 74348
rect 52237 74532 52293 74588
rect 52237 74452 52293 74508
rect 52237 74372 52293 74428
rect 52237 74292 52293 74348
rect 53638 74532 53694 74588
rect 53638 74452 53694 74508
rect 53638 74372 53694 74428
rect 53638 74292 53694 74348
rect 53806 74532 53862 74588
rect 53806 74452 53862 74508
rect 53806 74372 53862 74428
rect 53806 74292 53862 74348
rect 54550 74532 54606 74588
rect 54550 74452 54606 74508
rect 54550 74372 54606 74428
rect 54550 74292 54606 74348
rect 54940 74532 54996 74588
rect 54940 74452 54996 74508
rect 54940 74372 54996 74428
rect 54940 74292 54996 74348
rect 55656 74532 55712 74588
rect 55656 74452 55712 74508
rect 55656 74372 55712 74428
rect 55656 74292 55712 74348
rect 56234 74532 56290 74588
rect 56234 74452 56290 74508
rect 56234 74372 56290 74428
rect 56234 74292 56290 74348
rect 56679 74532 56735 74588
rect 56679 74452 56735 74508
rect 56679 74372 56735 74428
rect 56679 74292 56735 74348
rect 56983 74532 57039 74588
rect 56983 74452 57039 74508
rect 56983 74372 57039 74428
rect 56983 74292 57039 74348
rect 57825 74532 57881 74588
rect 57825 74452 57881 74508
rect 57825 74372 57881 74428
rect 57825 74292 57881 74348
rect 58465 74532 58521 74588
rect 58465 74452 58521 74508
rect 58465 74372 58521 74428
rect 58465 74292 58521 74348
rect 59048 74532 59104 74588
rect 59048 74452 59104 74508
rect 59048 74372 59104 74428
rect 59048 74292 59104 74348
rect 60326 74532 60382 74588
rect 60326 74452 60382 74508
rect 60326 74372 60382 74428
rect 60326 74292 60382 74348
rect 60484 74532 60540 74588
rect 60484 74452 60540 74508
rect 60484 74372 60540 74428
rect 60484 74292 60540 74348
rect 62528 74532 62584 74588
rect 62608 74532 62664 74588
rect 62528 74452 62584 74508
rect 62608 74452 62664 74508
rect 62528 74372 62584 74428
rect 62608 74372 62664 74428
rect 62528 74292 62584 74348
rect 62608 74292 62664 74348
rect 2184 72180 2240 72236
rect 2264 72180 2320 72236
rect 2184 72100 2240 72156
rect 2264 72100 2320 72156
rect 2184 72020 2240 72076
rect 2264 72020 2320 72076
rect 2184 71940 2240 71996
rect 2264 71940 2320 71996
rect 5393 72180 5449 72236
rect 5393 72100 5449 72156
rect 5393 72020 5449 72076
rect 5393 71940 5449 71996
rect 8283 72180 8339 72236
rect 8283 72100 8339 72156
rect 8283 72020 8339 72076
rect 8283 71940 8339 71996
rect 11173 72180 11229 72236
rect 11173 72100 11229 72156
rect 11173 72020 11229 72076
rect 11173 71940 11229 71996
rect 14063 72180 14119 72236
rect 14063 72100 14119 72156
rect 14063 72020 14119 72076
rect 14063 71940 14119 71996
rect 16953 72180 17009 72236
rect 16953 72100 17009 72156
rect 16953 72020 17009 72076
rect 16953 71940 17009 71996
rect 19843 72180 19899 72236
rect 19843 72100 19899 72156
rect 19843 72020 19899 72076
rect 19843 71940 19899 71996
rect 22733 72180 22789 72236
rect 22733 72100 22789 72156
rect 22733 72020 22789 72076
rect 22733 71940 22789 71996
rect 25623 72180 25679 72236
rect 25623 72100 25679 72156
rect 25623 72020 25679 72076
rect 25623 71940 25679 71996
rect 28513 72180 28569 72236
rect 28513 72100 28569 72156
rect 28513 72020 28569 72076
rect 28513 71940 28569 71996
rect 31403 72180 31459 72236
rect 31403 72100 31459 72156
rect 31403 72020 31459 72076
rect 31403 71940 31459 71996
rect 34293 72180 34349 72236
rect 34293 72100 34349 72156
rect 34293 72020 34349 72076
rect 34293 71940 34349 71996
rect 37183 72180 37239 72236
rect 37183 72100 37239 72156
rect 37183 72020 37239 72076
rect 37183 71940 37239 71996
rect 40073 72180 40129 72236
rect 40073 72100 40129 72156
rect 40073 72020 40129 72076
rect 40073 71940 40129 71996
rect 42963 72180 43019 72236
rect 42963 72100 43019 72156
rect 42963 72020 43019 72076
rect 42963 71940 43019 71996
rect 45853 72180 45909 72236
rect 45853 72100 45909 72156
rect 45853 72020 45909 72076
rect 45853 71940 45909 71996
rect 48800 72180 48856 72236
rect 48800 72100 48856 72156
rect 48800 72020 48856 72076
rect 48800 71940 48856 71996
rect 49662 72180 49718 72236
rect 49742 72180 49798 72236
rect 49662 72100 49718 72156
rect 49742 72100 49798 72156
rect 49662 72020 49718 72076
rect 49742 72020 49798 72076
rect 49662 71940 49718 71996
rect 49742 71940 49798 71996
rect 52956 72180 53012 72236
rect 52956 72100 53012 72156
rect 52956 72020 53012 72076
rect 52956 71940 53012 71996
rect 53114 72180 53170 72236
rect 53114 72100 53170 72156
rect 53114 72020 53170 72076
rect 53114 71940 53170 71996
rect 53470 72180 53526 72236
rect 53470 72100 53526 72156
rect 53470 72020 53526 72076
rect 53470 71940 53526 71996
rect 54788 72180 54844 72236
rect 54788 72100 54844 72156
rect 54788 72020 54844 72076
rect 54788 71940 54844 71996
rect 55381 72180 55437 72236
rect 55381 72100 55437 72156
rect 55381 72020 55437 72076
rect 55381 71940 55437 71996
rect 56527 72180 56583 72236
rect 56527 72100 56583 72156
rect 56527 72020 56583 72076
rect 56527 71940 56583 71996
rect 57963 72180 58019 72236
rect 58043 72180 58099 72236
rect 57963 72100 58019 72156
rect 58043 72100 58099 72156
rect 57963 72020 58019 72076
rect 58043 72020 58099 72076
rect 57963 71940 58019 71996
rect 58043 71940 58099 71996
rect 59206 72180 59262 72236
rect 59206 72100 59262 72156
rect 59206 72020 59262 72076
rect 59206 71940 59262 71996
rect 59364 72180 59420 72236
rect 59364 72100 59420 72156
rect 59364 72020 59420 72076
rect 59364 71940 59420 71996
rect 59672 72180 59728 72236
rect 59672 72100 59728 72156
rect 59672 72020 59728 72076
rect 59672 71940 59728 71996
rect 59818 72180 59874 72236
rect 59818 72100 59874 72156
rect 59818 72020 59874 72076
rect 59818 71940 59874 71996
rect 59954 72180 60010 72236
rect 60034 72180 60090 72236
rect 59954 72100 60010 72156
rect 60034 72100 60090 72156
rect 59954 72020 60010 72076
rect 60034 72020 60090 72076
rect 59954 71940 60010 71996
rect 60034 71940 60090 71996
rect 62326 72180 62382 72236
rect 62406 72180 62462 72236
rect 62326 72100 62382 72156
rect 62406 72100 62462 72156
rect 62326 72020 62382 72076
rect 62406 72020 62462 72076
rect 62326 71940 62382 71996
rect 62406 71940 62462 71996
rect 2044 64532 2100 64588
rect 2044 64452 2100 64508
rect 2044 64372 2100 64428
rect 2044 64292 2100 64348
rect 5540 64532 5596 64588
rect 5540 64452 5596 64508
rect 5540 64372 5596 64428
rect 5540 64292 5596 64348
rect 8430 64532 8486 64588
rect 8430 64452 8486 64508
rect 8430 64372 8486 64428
rect 8430 64292 8486 64348
rect 11320 64532 11376 64588
rect 11320 64452 11376 64508
rect 11320 64372 11376 64428
rect 11320 64292 11376 64348
rect 14210 64532 14266 64588
rect 14210 64452 14266 64508
rect 14210 64372 14266 64428
rect 14210 64292 14266 64348
rect 17100 64532 17156 64588
rect 17100 64452 17156 64508
rect 17100 64372 17156 64428
rect 17100 64292 17156 64348
rect 19990 64532 20046 64588
rect 19990 64452 20046 64508
rect 19990 64372 20046 64428
rect 19990 64292 20046 64348
rect 22880 64532 22936 64588
rect 22880 64452 22936 64508
rect 22880 64372 22936 64428
rect 22880 64292 22936 64348
rect 25770 64532 25826 64588
rect 25770 64452 25826 64508
rect 25770 64372 25826 64428
rect 25770 64292 25826 64348
rect 28660 64532 28716 64588
rect 28660 64452 28716 64508
rect 28660 64372 28716 64428
rect 28660 64292 28716 64348
rect 31550 64532 31606 64588
rect 31550 64452 31606 64508
rect 31550 64372 31606 64428
rect 31550 64292 31606 64348
rect 34440 64532 34496 64588
rect 34440 64452 34496 64508
rect 34440 64372 34496 64428
rect 34440 64292 34496 64348
rect 37330 64532 37386 64588
rect 37330 64452 37386 64508
rect 37330 64372 37386 64428
rect 37330 64292 37386 64348
rect 40220 64532 40276 64588
rect 40220 64452 40276 64508
rect 40220 64372 40276 64428
rect 40220 64292 40276 64348
rect 43110 64532 43166 64588
rect 43110 64452 43166 64508
rect 43110 64372 43166 64428
rect 43110 64292 43166 64348
rect 46000 64532 46056 64588
rect 46000 64452 46056 64508
rect 46000 64372 46056 64428
rect 46000 64292 46056 64348
rect 49008 64532 49064 64588
rect 49008 64452 49064 64508
rect 49008 64372 49064 64428
rect 49008 64292 49064 64348
rect 52237 64532 52293 64588
rect 52237 64452 52293 64508
rect 52237 64372 52293 64428
rect 52237 64292 52293 64348
rect 53638 64532 53694 64588
rect 53638 64452 53694 64508
rect 53638 64372 53694 64428
rect 53638 64292 53694 64348
rect 53806 64532 53862 64588
rect 53806 64452 53862 64508
rect 53806 64372 53862 64428
rect 53806 64292 53862 64348
rect 54550 64532 54606 64588
rect 54550 64452 54606 64508
rect 54550 64372 54606 64428
rect 54550 64292 54606 64348
rect 54940 64532 54996 64588
rect 54940 64452 54996 64508
rect 54940 64372 54996 64428
rect 54940 64292 54996 64348
rect 55656 64532 55712 64588
rect 55656 64452 55712 64508
rect 55656 64372 55712 64428
rect 55656 64292 55712 64348
rect 56234 64532 56290 64588
rect 56234 64452 56290 64508
rect 56234 64372 56290 64428
rect 56234 64292 56290 64348
rect 56679 64532 56735 64588
rect 56679 64452 56735 64508
rect 56679 64372 56735 64428
rect 56679 64292 56735 64348
rect 56983 64532 57039 64588
rect 56983 64452 57039 64508
rect 56983 64372 57039 64428
rect 56983 64292 57039 64348
rect 57825 64532 57881 64588
rect 57825 64452 57881 64508
rect 57825 64372 57881 64428
rect 57825 64292 57881 64348
rect 58465 64532 58521 64588
rect 58465 64452 58521 64508
rect 58465 64372 58521 64428
rect 58465 64292 58521 64348
rect 59048 64532 59104 64588
rect 59048 64452 59104 64508
rect 59048 64372 59104 64428
rect 59048 64292 59104 64348
rect 60326 64532 60382 64588
rect 60326 64452 60382 64508
rect 60326 64372 60382 64428
rect 60326 64292 60382 64348
rect 60484 64532 60540 64588
rect 60484 64452 60540 64508
rect 60484 64372 60540 64428
rect 60484 64292 60540 64348
rect 62528 64532 62584 64588
rect 62608 64532 62664 64588
rect 62528 64452 62584 64508
rect 62608 64452 62664 64508
rect 62528 64372 62584 64428
rect 62608 64372 62664 64428
rect 62528 64292 62584 64348
rect 62608 64292 62664 64348
rect 2184 62180 2240 62236
rect 2264 62180 2320 62236
rect 2184 62100 2240 62156
rect 2264 62100 2320 62156
rect 2184 62020 2240 62076
rect 2264 62020 2320 62076
rect 2184 61940 2240 61996
rect 2264 61940 2320 61996
rect 5393 62180 5449 62236
rect 5393 62100 5449 62156
rect 5393 62020 5449 62076
rect 5393 61940 5449 61996
rect 8283 62180 8339 62236
rect 8283 62100 8339 62156
rect 8283 62020 8339 62076
rect 8283 61940 8339 61996
rect 11173 62180 11229 62236
rect 11173 62100 11229 62156
rect 11173 62020 11229 62076
rect 11173 61940 11229 61996
rect 14063 62180 14119 62236
rect 14063 62100 14119 62156
rect 14063 62020 14119 62076
rect 14063 61940 14119 61996
rect 16953 62180 17009 62236
rect 16953 62100 17009 62156
rect 16953 62020 17009 62076
rect 16953 61940 17009 61996
rect 19843 62180 19899 62236
rect 19843 62100 19899 62156
rect 19843 62020 19899 62076
rect 19843 61940 19899 61996
rect 22733 62180 22789 62236
rect 22733 62100 22789 62156
rect 22733 62020 22789 62076
rect 22733 61940 22789 61996
rect 25623 62180 25679 62236
rect 25623 62100 25679 62156
rect 25623 62020 25679 62076
rect 25623 61940 25679 61996
rect 28513 62180 28569 62236
rect 28513 62100 28569 62156
rect 28513 62020 28569 62076
rect 28513 61940 28569 61996
rect 31403 62180 31459 62236
rect 31403 62100 31459 62156
rect 31403 62020 31459 62076
rect 31403 61940 31459 61996
rect 34293 62180 34349 62236
rect 34293 62100 34349 62156
rect 34293 62020 34349 62076
rect 34293 61940 34349 61996
rect 37183 62180 37239 62236
rect 37183 62100 37239 62156
rect 37183 62020 37239 62076
rect 37183 61940 37239 61996
rect 40073 62180 40129 62236
rect 40073 62100 40129 62156
rect 40073 62020 40129 62076
rect 40073 61940 40129 61996
rect 42963 62180 43019 62236
rect 42963 62100 43019 62156
rect 42963 62020 43019 62076
rect 42963 61940 43019 61996
rect 45853 62180 45909 62236
rect 45853 62100 45909 62156
rect 45853 62020 45909 62076
rect 45853 61940 45909 61996
rect 48800 62180 48856 62236
rect 48800 62100 48856 62156
rect 48800 62020 48856 62076
rect 48800 61940 48856 61996
rect 49662 62180 49718 62236
rect 49742 62180 49798 62236
rect 49662 62100 49718 62156
rect 49742 62100 49798 62156
rect 49662 62020 49718 62076
rect 49742 62020 49798 62076
rect 49662 61940 49718 61996
rect 49742 61940 49798 61996
rect 52956 62180 53012 62236
rect 52956 62100 53012 62156
rect 52956 62020 53012 62076
rect 52956 61940 53012 61996
rect 53114 62180 53170 62236
rect 53114 62100 53170 62156
rect 53114 62020 53170 62076
rect 53114 61940 53170 61996
rect 53470 62180 53526 62236
rect 53470 62100 53526 62156
rect 53470 62020 53526 62076
rect 53470 61940 53526 61996
rect 54788 62180 54844 62236
rect 54788 62100 54844 62156
rect 54788 62020 54844 62076
rect 54788 61940 54844 61996
rect 55381 62180 55437 62236
rect 55381 62100 55437 62156
rect 55381 62020 55437 62076
rect 55381 61940 55437 61996
rect 56527 62180 56583 62236
rect 56527 62100 56583 62156
rect 56527 62020 56583 62076
rect 56527 61940 56583 61996
rect 57963 62180 58019 62236
rect 58043 62180 58099 62236
rect 57963 62100 58019 62156
rect 58043 62100 58099 62156
rect 57963 62020 58019 62076
rect 58043 62020 58099 62076
rect 57963 61940 58019 61996
rect 58043 61940 58099 61996
rect 59206 62180 59262 62236
rect 59206 62100 59262 62156
rect 59206 62020 59262 62076
rect 59206 61940 59262 61996
rect 59364 62180 59420 62236
rect 59364 62100 59420 62156
rect 59364 62020 59420 62076
rect 59364 61940 59420 61996
rect 59672 62180 59728 62236
rect 59672 62100 59728 62156
rect 59672 62020 59728 62076
rect 59672 61940 59728 61996
rect 59818 62180 59874 62236
rect 59818 62100 59874 62156
rect 59818 62020 59874 62076
rect 59818 61940 59874 61996
rect 59954 62180 60010 62236
rect 60034 62180 60090 62236
rect 59954 62100 60010 62156
rect 60034 62100 60090 62156
rect 59954 62020 60010 62076
rect 60034 62020 60090 62076
rect 59954 61940 60010 61996
rect 60034 61940 60090 61996
rect 62326 62180 62382 62236
rect 62406 62180 62462 62236
rect 62326 62100 62382 62156
rect 62406 62100 62462 62156
rect 62326 62020 62382 62076
rect 62406 62020 62462 62076
rect 62326 61940 62382 61996
rect 62406 61940 62462 61996
rect 2044 54532 2100 54588
rect 2044 54452 2100 54508
rect 2044 54372 2100 54428
rect 2044 54292 2100 54348
rect 5540 54532 5596 54588
rect 5540 54452 5596 54508
rect 5540 54372 5596 54428
rect 5540 54292 5596 54348
rect 8430 54532 8486 54588
rect 8430 54452 8486 54508
rect 8430 54372 8486 54428
rect 8430 54292 8486 54348
rect 11320 54532 11376 54588
rect 11320 54452 11376 54508
rect 11320 54372 11376 54428
rect 11320 54292 11376 54348
rect 14210 54532 14266 54588
rect 14210 54452 14266 54508
rect 14210 54372 14266 54428
rect 14210 54292 14266 54348
rect 17100 54532 17156 54588
rect 17100 54452 17156 54508
rect 17100 54372 17156 54428
rect 17100 54292 17156 54348
rect 19990 54532 20046 54588
rect 19990 54452 20046 54508
rect 19990 54372 20046 54428
rect 19990 54292 20046 54348
rect 22880 54532 22936 54588
rect 22880 54452 22936 54508
rect 22880 54372 22936 54428
rect 22880 54292 22936 54348
rect 25770 54532 25826 54588
rect 25770 54452 25826 54508
rect 25770 54372 25826 54428
rect 25770 54292 25826 54348
rect 28660 54532 28716 54588
rect 28660 54452 28716 54508
rect 28660 54372 28716 54428
rect 28660 54292 28716 54348
rect 31550 54532 31606 54588
rect 31550 54452 31606 54508
rect 31550 54372 31606 54428
rect 31550 54292 31606 54348
rect 34440 54532 34496 54588
rect 34440 54452 34496 54508
rect 34440 54372 34496 54428
rect 34440 54292 34496 54348
rect 37330 54532 37386 54588
rect 37330 54452 37386 54508
rect 37330 54372 37386 54428
rect 37330 54292 37386 54348
rect 40220 54532 40276 54588
rect 40220 54452 40276 54508
rect 40220 54372 40276 54428
rect 40220 54292 40276 54348
rect 43110 54532 43166 54588
rect 43110 54452 43166 54508
rect 43110 54372 43166 54428
rect 43110 54292 43166 54348
rect 46000 54532 46056 54588
rect 46000 54452 46056 54508
rect 46000 54372 46056 54428
rect 46000 54292 46056 54348
rect 49008 54532 49064 54588
rect 49008 54452 49064 54508
rect 49008 54372 49064 54428
rect 49008 54292 49064 54348
rect 52237 54532 52293 54588
rect 52237 54452 52293 54508
rect 52237 54372 52293 54428
rect 52237 54292 52293 54348
rect 53638 54532 53694 54588
rect 53638 54452 53694 54508
rect 53638 54372 53694 54428
rect 53638 54292 53694 54348
rect 53806 54532 53862 54588
rect 53806 54452 53862 54508
rect 53806 54372 53862 54428
rect 53806 54292 53862 54348
rect 54550 54532 54606 54588
rect 54550 54452 54606 54508
rect 54550 54372 54606 54428
rect 54550 54292 54606 54348
rect 54940 54532 54996 54588
rect 54940 54452 54996 54508
rect 54940 54372 54996 54428
rect 54940 54292 54996 54348
rect 55656 54532 55712 54588
rect 55656 54452 55712 54508
rect 55656 54372 55712 54428
rect 55656 54292 55712 54348
rect 56234 54532 56290 54588
rect 56234 54452 56290 54508
rect 56234 54372 56290 54428
rect 56234 54292 56290 54348
rect 56679 54532 56735 54588
rect 56679 54452 56735 54508
rect 56679 54372 56735 54428
rect 56679 54292 56735 54348
rect 56983 54532 57039 54588
rect 56983 54452 57039 54508
rect 56983 54372 57039 54428
rect 56983 54292 57039 54348
rect 57825 54532 57881 54588
rect 57825 54452 57881 54508
rect 57825 54372 57881 54428
rect 57825 54292 57881 54348
rect 58465 54532 58521 54588
rect 58465 54452 58521 54508
rect 58465 54372 58521 54428
rect 58465 54292 58521 54348
rect 59048 54532 59104 54588
rect 59048 54452 59104 54508
rect 59048 54372 59104 54428
rect 59048 54292 59104 54348
rect 60326 54532 60382 54588
rect 60326 54452 60382 54508
rect 60326 54372 60382 54428
rect 60326 54292 60382 54348
rect 60484 54532 60540 54588
rect 60484 54452 60540 54508
rect 60484 54372 60540 54428
rect 60484 54292 60540 54348
rect 62528 54532 62584 54588
rect 62608 54532 62664 54588
rect 62528 54452 62584 54508
rect 62608 54452 62664 54508
rect 62528 54372 62584 54428
rect 62608 54372 62664 54428
rect 62528 54292 62584 54348
rect 62608 54292 62664 54348
rect 2184 52180 2240 52236
rect 2264 52180 2320 52236
rect 2184 52100 2240 52156
rect 2264 52100 2320 52156
rect 2184 52020 2240 52076
rect 2264 52020 2320 52076
rect 2184 51940 2240 51996
rect 2264 51940 2320 51996
rect 5393 52180 5449 52236
rect 5393 52100 5449 52156
rect 5393 52020 5449 52076
rect 5393 51940 5449 51996
rect 8283 52180 8339 52236
rect 8283 52100 8339 52156
rect 8283 52020 8339 52076
rect 8283 51940 8339 51996
rect 11173 52180 11229 52236
rect 11173 52100 11229 52156
rect 11173 52020 11229 52076
rect 11173 51940 11229 51996
rect 14063 52180 14119 52236
rect 14063 52100 14119 52156
rect 14063 52020 14119 52076
rect 14063 51940 14119 51996
rect 16953 52180 17009 52236
rect 16953 52100 17009 52156
rect 16953 52020 17009 52076
rect 16953 51940 17009 51996
rect 19843 52180 19899 52236
rect 19843 52100 19899 52156
rect 19843 52020 19899 52076
rect 19843 51940 19899 51996
rect 22733 52180 22789 52236
rect 22733 52100 22789 52156
rect 22733 52020 22789 52076
rect 22733 51940 22789 51996
rect 25623 52180 25679 52236
rect 25623 52100 25679 52156
rect 25623 52020 25679 52076
rect 25623 51940 25679 51996
rect 28513 52180 28569 52236
rect 28513 52100 28569 52156
rect 28513 52020 28569 52076
rect 28513 51940 28569 51996
rect 31403 52180 31459 52236
rect 31403 52100 31459 52156
rect 31403 52020 31459 52076
rect 31403 51940 31459 51996
rect 34293 52180 34349 52236
rect 34293 52100 34349 52156
rect 34293 52020 34349 52076
rect 34293 51940 34349 51996
rect 37183 52180 37239 52236
rect 37183 52100 37239 52156
rect 37183 52020 37239 52076
rect 37183 51940 37239 51996
rect 40073 52180 40129 52236
rect 40073 52100 40129 52156
rect 40073 52020 40129 52076
rect 40073 51940 40129 51996
rect 42963 52180 43019 52236
rect 42963 52100 43019 52156
rect 42963 52020 43019 52076
rect 42963 51940 43019 51996
rect 45853 52180 45909 52236
rect 45853 52100 45909 52156
rect 45853 52020 45909 52076
rect 45853 51940 45909 51996
rect 48800 52180 48856 52236
rect 48800 52100 48856 52156
rect 48800 52020 48856 52076
rect 48800 51940 48856 51996
rect 49662 52180 49718 52236
rect 49742 52180 49798 52236
rect 49662 52100 49718 52156
rect 49742 52100 49798 52156
rect 49662 52020 49718 52076
rect 49742 52020 49798 52076
rect 49662 51940 49718 51996
rect 49742 51940 49798 51996
rect 52956 52180 53012 52236
rect 52956 52100 53012 52156
rect 52956 52020 53012 52076
rect 52956 51940 53012 51996
rect 53114 52180 53170 52236
rect 53114 52100 53170 52156
rect 53114 52020 53170 52076
rect 53114 51940 53170 51996
rect 53470 52180 53526 52236
rect 53470 52100 53526 52156
rect 53470 52020 53526 52076
rect 53470 51940 53526 51996
rect 54788 52180 54844 52236
rect 54788 52100 54844 52156
rect 54788 52020 54844 52076
rect 54788 51940 54844 51996
rect 55381 52180 55437 52236
rect 55381 52100 55437 52156
rect 55381 52020 55437 52076
rect 55381 51940 55437 51996
rect 56527 52180 56583 52236
rect 56527 52100 56583 52156
rect 56527 52020 56583 52076
rect 56527 51940 56583 51996
rect 57963 52180 58019 52236
rect 58043 52180 58099 52236
rect 57963 52100 58019 52156
rect 58043 52100 58099 52156
rect 57963 52020 58019 52076
rect 58043 52020 58099 52076
rect 57963 51940 58019 51996
rect 58043 51940 58099 51996
rect 59206 52180 59262 52236
rect 59206 52100 59262 52156
rect 59206 52020 59262 52076
rect 59206 51940 59262 51996
rect 59364 52180 59420 52236
rect 59364 52100 59420 52156
rect 59364 52020 59420 52076
rect 59364 51940 59420 51996
rect 59672 52180 59728 52236
rect 59672 52100 59728 52156
rect 59672 52020 59728 52076
rect 59672 51940 59728 51996
rect 59818 52180 59874 52236
rect 59818 52100 59874 52156
rect 59818 52020 59874 52076
rect 59818 51940 59874 51996
rect 59954 52180 60010 52236
rect 60034 52180 60090 52236
rect 59954 52100 60010 52156
rect 60034 52100 60090 52156
rect 59954 52020 60010 52076
rect 60034 52020 60090 52076
rect 59954 51940 60010 51996
rect 60034 51940 60090 51996
rect 62326 52180 62382 52236
rect 62406 52180 62462 52236
rect 62326 52100 62382 52156
rect 62406 52100 62462 52156
rect 62326 52020 62382 52076
rect 62406 52020 62462 52076
rect 62326 51940 62382 51996
rect 62406 51940 62462 51996
rect 2044 44532 2100 44588
rect 2044 44452 2100 44508
rect 2044 44372 2100 44428
rect 2044 44292 2100 44348
rect 5540 44532 5596 44588
rect 5540 44452 5596 44508
rect 5540 44372 5596 44428
rect 5540 44292 5596 44348
rect 8430 44532 8486 44588
rect 8430 44452 8486 44508
rect 8430 44372 8486 44428
rect 8430 44292 8486 44348
rect 11320 44532 11376 44588
rect 11320 44452 11376 44508
rect 11320 44372 11376 44428
rect 11320 44292 11376 44348
rect 14210 44532 14266 44588
rect 14210 44452 14266 44508
rect 14210 44372 14266 44428
rect 14210 44292 14266 44348
rect 17100 44532 17156 44588
rect 17100 44452 17156 44508
rect 17100 44372 17156 44428
rect 17100 44292 17156 44348
rect 19990 44532 20046 44588
rect 19990 44452 20046 44508
rect 19990 44372 20046 44428
rect 19990 44292 20046 44348
rect 22880 44532 22936 44588
rect 22880 44452 22936 44508
rect 22880 44372 22936 44428
rect 22880 44292 22936 44348
rect 25770 44532 25826 44588
rect 25770 44452 25826 44508
rect 25770 44372 25826 44428
rect 25770 44292 25826 44348
rect 28660 44532 28716 44588
rect 28660 44452 28716 44508
rect 28660 44372 28716 44428
rect 28660 44292 28716 44348
rect 31550 44532 31606 44588
rect 31550 44452 31606 44508
rect 31550 44372 31606 44428
rect 31550 44292 31606 44348
rect 34440 44532 34496 44588
rect 34440 44452 34496 44508
rect 34440 44372 34496 44428
rect 34440 44292 34496 44348
rect 37330 44532 37386 44588
rect 37330 44452 37386 44508
rect 37330 44372 37386 44428
rect 37330 44292 37386 44348
rect 40220 44532 40276 44588
rect 40220 44452 40276 44508
rect 40220 44372 40276 44428
rect 40220 44292 40276 44348
rect 43110 44532 43166 44588
rect 43110 44452 43166 44508
rect 43110 44372 43166 44428
rect 43110 44292 43166 44348
rect 46000 44532 46056 44588
rect 46000 44452 46056 44508
rect 46000 44372 46056 44428
rect 46000 44292 46056 44348
rect 52237 44532 52293 44588
rect 52237 44452 52293 44508
rect 52237 44372 52293 44428
rect 52237 44292 52293 44348
rect 53638 44532 53694 44588
rect 53638 44452 53694 44508
rect 53638 44372 53694 44428
rect 53638 44292 53694 44348
rect 54550 44532 54606 44588
rect 54550 44452 54606 44508
rect 54550 44372 54606 44428
rect 54550 44292 54606 44348
rect 54940 44532 54996 44588
rect 54940 44452 54996 44508
rect 54940 44372 54996 44428
rect 54940 44292 54996 44348
rect 55656 44532 55712 44588
rect 55656 44452 55712 44508
rect 55656 44372 55712 44428
rect 55656 44292 55712 44348
rect 56234 44532 56290 44588
rect 56234 44452 56290 44508
rect 56234 44372 56290 44428
rect 56234 44292 56290 44348
rect 56679 44532 56735 44588
rect 56679 44452 56735 44508
rect 56679 44372 56735 44428
rect 56679 44292 56735 44348
rect 56983 44532 57039 44588
rect 56983 44452 57039 44508
rect 56983 44372 57039 44428
rect 56983 44292 57039 44348
rect 57825 44532 57881 44588
rect 57825 44452 57881 44508
rect 57825 44372 57881 44428
rect 57825 44292 57881 44348
rect 58349 44532 58405 44588
rect 58349 44452 58405 44508
rect 58349 44372 58405 44428
rect 58349 44292 58405 44348
rect 59048 44532 59104 44588
rect 59048 44452 59104 44508
rect 59048 44372 59104 44428
rect 59048 44292 59104 44348
rect 60326 44532 60382 44588
rect 60326 44452 60382 44508
rect 60326 44372 60382 44428
rect 60326 44292 60382 44348
rect 60484 44532 60540 44588
rect 60484 44452 60540 44508
rect 60484 44372 60540 44428
rect 60484 44292 60540 44348
rect 62528 44532 62584 44588
rect 62608 44532 62664 44588
rect 62528 44452 62584 44508
rect 62608 44452 62664 44508
rect 62528 44372 62584 44428
rect 62608 44372 62664 44428
rect 62528 44292 62584 44348
rect 62608 44292 62664 44348
rect 2184 42180 2240 42236
rect 2264 42180 2320 42236
rect 2184 42100 2240 42156
rect 2264 42100 2320 42156
rect 2184 42020 2240 42076
rect 2264 42020 2320 42076
rect 2184 41940 2240 41996
rect 2264 41940 2320 41996
rect 5393 42180 5449 42236
rect 5393 42100 5449 42156
rect 5393 42020 5449 42076
rect 5393 41940 5449 41996
rect 8283 42180 8339 42236
rect 8283 42100 8339 42156
rect 8283 42020 8339 42076
rect 8283 41940 8339 41996
rect 11173 42180 11229 42236
rect 11173 42100 11229 42156
rect 11173 42020 11229 42076
rect 11173 41940 11229 41996
rect 14063 42180 14119 42236
rect 14063 42100 14119 42156
rect 14063 42020 14119 42076
rect 14063 41940 14119 41996
rect 16953 42180 17009 42236
rect 16953 42100 17009 42156
rect 16953 42020 17009 42076
rect 16953 41940 17009 41996
rect 19843 42180 19899 42236
rect 19843 42100 19899 42156
rect 19843 42020 19899 42076
rect 19843 41940 19899 41996
rect 22733 42180 22789 42236
rect 22733 42100 22789 42156
rect 22733 42020 22789 42076
rect 22733 41940 22789 41996
rect 25623 42180 25679 42236
rect 25623 42100 25679 42156
rect 25623 42020 25679 42076
rect 25623 41940 25679 41996
rect 28513 42180 28569 42236
rect 28513 42100 28569 42156
rect 28513 42020 28569 42076
rect 28513 41940 28569 41996
rect 31403 42180 31459 42236
rect 31403 42100 31459 42156
rect 31403 42020 31459 42076
rect 31403 41940 31459 41996
rect 34293 42180 34349 42236
rect 34293 42100 34349 42156
rect 34293 42020 34349 42076
rect 34293 41940 34349 41996
rect 37183 42180 37239 42236
rect 37183 42100 37239 42156
rect 37183 42020 37239 42076
rect 37183 41940 37239 41996
rect 40073 42180 40129 42236
rect 40073 42100 40129 42156
rect 40073 42020 40129 42076
rect 40073 41940 40129 41996
rect 42963 42180 43019 42236
rect 42963 42100 43019 42156
rect 42963 42020 43019 42076
rect 42963 41940 43019 41996
rect 45853 42180 45909 42236
rect 45853 42100 45909 42156
rect 45853 42020 45909 42076
rect 45853 41940 45909 41996
rect 48800 42180 48856 42236
rect 48800 42100 48856 42156
rect 48800 42020 48856 42076
rect 48800 41940 48856 41996
rect 49662 42180 49718 42236
rect 49742 42180 49798 42236
rect 49662 42100 49718 42156
rect 49742 42100 49798 42156
rect 49662 42020 49718 42076
rect 49742 42020 49798 42076
rect 49662 41940 49718 41996
rect 49742 41940 49798 41996
rect 52956 42180 53012 42236
rect 52956 42100 53012 42156
rect 52956 42020 53012 42076
rect 52956 41940 53012 41996
rect 53114 42180 53170 42236
rect 53114 42100 53170 42156
rect 53114 42020 53170 42076
rect 53114 41940 53170 41996
rect 53470 42180 53526 42236
rect 53470 42100 53526 42156
rect 53470 42020 53526 42076
rect 53470 41940 53526 41996
rect 54788 42180 54844 42236
rect 54788 42100 54844 42156
rect 54788 42020 54844 42076
rect 54788 41940 54844 41996
rect 55381 42180 55437 42236
rect 55381 42100 55437 42156
rect 55381 42020 55437 42076
rect 55381 41940 55437 41996
rect 56527 42180 56583 42236
rect 56527 42100 56583 42156
rect 56527 42020 56583 42076
rect 56527 41940 56583 41996
rect 57963 42180 58019 42236
rect 58043 42180 58099 42236
rect 57963 42100 58019 42156
rect 58043 42100 58099 42156
rect 57963 42020 58019 42076
rect 58043 42020 58099 42076
rect 57963 41940 58019 41996
rect 58043 41940 58099 41996
rect 59206 42180 59262 42236
rect 59206 42100 59262 42156
rect 59206 42020 59262 42076
rect 59206 41940 59262 41996
rect 59364 42180 59420 42236
rect 59364 42100 59420 42156
rect 59364 42020 59420 42076
rect 59364 41940 59420 41996
rect 59672 42180 59728 42236
rect 59672 42100 59728 42156
rect 59672 42020 59728 42076
rect 59672 41940 59728 41996
rect 59818 42180 59874 42236
rect 59818 42100 59874 42156
rect 59818 42020 59874 42076
rect 59818 41940 59874 41996
rect 59954 42180 60010 42236
rect 60034 42180 60090 42236
rect 59954 42100 60010 42156
rect 60034 42100 60090 42156
rect 59954 42020 60010 42076
rect 60034 42020 60090 42076
rect 59954 41940 60010 41996
rect 60034 41940 60090 41996
rect 62326 42180 62382 42236
rect 62406 42180 62462 42236
rect 62326 42100 62382 42156
rect 62406 42100 62462 42156
rect 62326 42020 62382 42076
rect 62406 42020 62462 42076
rect 62326 41940 62382 41996
rect 62406 41940 62462 41996
rect 2044 34532 2100 34588
rect 2044 34452 2100 34508
rect 2044 34372 2100 34428
rect 2044 34292 2100 34348
rect 5540 34532 5596 34588
rect 5540 34452 5596 34508
rect 5540 34372 5596 34428
rect 5540 34292 5596 34348
rect 8430 34532 8486 34588
rect 8430 34452 8486 34508
rect 8430 34372 8486 34428
rect 8430 34292 8486 34348
rect 11320 34532 11376 34588
rect 11320 34452 11376 34508
rect 11320 34372 11376 34428
rect 11320 34292 11376 34348
rect 14210 34532 14266 34588
rect 14210 34452 14266 34508
rect 14210 34372 14266 34428
rect 14210 34292 14266 34348
rect 17100 34532 17156 34588
rect 17100 34452 17156 34508
rect 17100 34372 17156 34428
rect 17100 34292 17156 34348
rect 19990 34532 20046 34588
rect 19990 34452 20046 34508
rect 19990 34372 20046 34428
rect 19990 34292 20046 34348
rect 22880 34532 22936 34588
rect 22880 34452 22936 34508
rect 22880 34372 22936 34428
rect 22880 34292 22936 34348
rect 25770 34532 25826 34588
rect 25770 34452 25826 34508
rect 25770 34372 25826 34428
rect 25770 34292 25826 34348
rect 28660 34532 28716 34588
rect 28660 34452 28716 34508
rect 28660 34372 28716 34428
rect 28660 34292 28716 34348
rect 31550 34532 31606 34588
rect 31550 34452 31606 34508
rect 31550 34372 31606 34428
rect 31550 34292 31606 34348
rect 34440 34532 34496 34588
rect 34440 34452 34496 34508
rect 34440 34372 34496 34428
rect 34440 34292 34496 34348
rect 37330 34532 37386 34588
rect 37330 34452 37386 34508
rect 37330 34372 37386 34428
rect 37330 34292 37386 34348
rect 40220 34532 40276 34588
rect 40220 34452 40276 34508
rect 40220 34372 40276 34428
rect 40220 34292 40276 34348
rect 43110 34532 43166 34588
rect 43110 34452 43166 34508
rect 43110 34372 43166 34428
rect 43110 34292 43166 34348
rect 46000 34532 46056 34588
rect 46000 34452 46056 34508
rect 46000 34372 46056 34428
rect 46000 34292 46056 34348
rect 49008 34532 49064 34588
rect 49008 34452 49064 34508
rect 49008 34372 49064 34428
rect 49008 34292 49064 34348
rect 52237 34532 52293 34588
rect 52237 34452 52293 34508
rect 52237 34372 52293 34428
rect 52237 34292 52293 34348
rect 53638 34532 53694 34588
rect 53638 34452 53694 34508
rect 53638 34372 53694 34428
rect 53638 34292 53694 34348
rect 53806 34532 53862 34588
rect 53806 34452 53862 34508
rect 53806 34372 53862 34428
rect 53806 34292 53862 34348
rect 54550 34532 54606 34588
rect 54550 34452 54606 34508
rect 54550 34372 54606 34428
rect 54550 34292 54606 34348
rect 54940 34532 54996 34588
rect 54940 34452 54996 34508
rect 54940 34372 54996 34428
rect 54940 34292 54996 34348
rect 55656 34532 55712 34588
rect 55656 34452 55712 34508
rect 55656 34372 55712 34428
rect 55656 34292 55712 34348
rect 56234 34532 56290 34588
rect 56234 34452 56290 34508
rect 56234 34372 56290 34428
rect 56234 34292 56290 34348
rect 56679 34532 56735 34588
rect 56679 34452 56735 34508
rect 56679 34372 56735 34428
rect 56679 34292 56735 34348
rect 56983 34532 57039 34588
rect 56983 34452 57039 34508
rect 56983 34372 57039 34428
rect 56983 34292 57039 34348
rect 57825 34532 57881 34588
rect 57825 34452 57881 34508
rect 57825 34372 57881 34428
rect 57825 34292 57881 34348
rect 58465 34532 58521 34588
rect 58465 34452 58521 34508
rect 58465 34372 58521 34428
rect 58465 34292 58521 34348
rect 59048 34532 59104 34588
rect 59048 34452 59104 34508
rect 59048 34372 59104 34428
rect 59048 34292 59104 34348
rect 60326 34532 60382 34588
rect 60326 34452 60382 34508
rect 60326 34372 60382 34428
rect 60326 34292 60382 34348
rect 60484 34532 60540 34588
rect 60484 34452 60540 34508
rect 60484 34372 60540 34428
rect 60484 34292 60540 34348
rect 62528 34532 62584 34588
rect 62608 34532 62664 34588
rect 62528 34452 62584 34508
rect 62608 34452 62664 34508
rect 62528 34372 62584 34428
rect 62608 34372 62664 34428
rect 62528 34292 62584 34348
rect 62608 34292 62664 34348
rect 2184 32180 2240 32236
rect 2264 32180 2320 32236
rect 2184 32100 2240 32156
rect 2264 32100 2320 32156
rect 2184 32020 2240 32076
rect 2264 32020 2320 32076
rect 2184 31940 2240 31996
rect 2264 31940 2320 31996
rect 5393 32180 5449 32236
rect 5393 32100 5449 32156
rect 5393 32020 5449 32076
rect 5393 31940 5449 31996
rect 8283 32180 8339 32236
rect 8283 32100 8339 32156
rect 8283 32020 8339 32076
rect 8283 31940 8339 31996
rect 11173 32180 11229 32236
rect 11173 32100 11229 32156
rect 11173 32020 11229 32076
rect 11173 31940 11229 31996
rect 14063 32180 14119 32236
rect 14063 32100 14119 32156
rect 14063 32020 14119 32076
rect 14063 31940 14119 31996
rect 16953 32180 17009 32236
rect 16953 32100 17009 32156
rect 16953 32020 17009 32076
rect 16953 31940 17009 31996
rect 19843 32180 19899 32236
rect 19843 32100 19899 32156
rect 19843 32020 19899 32076
rect 19843 31940 19899 31996
rect 22733 32180 22789 32236
rect 22733 32100 22789 32156
rect 22733 32020 22789 32076
rect 22733 31940 22789 31996
rect 25623 32180 25679 32236
rect 25623 32100 25679 32156
rect 25623 32020 25679 32076
rect 25623 31940 25679 31996
rect 28513 32180 28569 32236
rect 28513 32100 28569 32156
rect 28513 32020 28569 32076
rect 28513 31940 28569 31996
rect 31403 32180 31459 32236
rect 31403 32100 31459 32156
rect 31403 32020 31459 32076
rect 31403 31940 31459 31996
rect 34293 32180 34349 32236
rect 34293 32100 34349 32156
rect 34293 32020 34349 32076
rect 34293 31940 34349 31996
rect 37183 32180 37239 32236
rect 37183 32100 37239 32156
rect 37183 32020 37239 32076
rect 37183 31940 37239 31996
rect 40073 32180 40129 32236
rect 40073 32100 40129 32156
rect 40073 32020 40129 32076
rect 40073 31940 40129 31996
rect 42963 32180 43019 32236
rect 42963 32100 43019 32156
rect 42963 32020 43019 32076
rect 42963 31940 43019 31996
rect 45853 32180 45909 32236
rect 45853 32100 45909 32156
rect 45853 32020 45909 32076
rect 45853 31940 45909 31996
rect 48800 32180 48856 32236
rect 48800 32100 48856 32156
rect 48800 32020 48856 32076
rect 48800 31940 48856 31996
rect 49662 32180 49718 32236
rect 49742 32180 49798 32236
rect 49662 32100 49718 32156
rect 49742 32100 49798 32156
rect 49662 32020 49718 32076
rect 49742 32020 49798 32076
rect 49662 31940 49718 31996
rect 49742 31940 49798 31996
rect 52956 32180 53012 32236
rect 52956 32100 53012 32156
rect 52956 32020 53012 32076
rect 52956 31940 53012 31996
rect 53114 32180 53170 32236
rect 53114 32100 53170 32156
rect 53114 32020 53170 32076
rect 53114 31940 53170 31996
rect 53470 32180 53526 32236
rect 53470 32100 53526 32156
rect 53470 32020 53526 32076
rect 53470 31940 53526 31996
rect 54788 32180 54844 32236
rect 54788 32100 54844 32156
rect 54788 32020 54844 32076
rect 54788 31940 54844 31996
rect 55381 32180 55437 32236
rect 55381 32100 55437 32156
rect 55381 32020 55437 32076
rect 55381 31940 55437 31996
rect 56527 32180 56583 32236
rect 56527 32100 56583 32156
rect 56527 32020 56583 32076
rect 56527 31940 56583 31996
rect 57963 32180 58019 32236
rect 58043 32180 58099 32236
rect 57963 32100 58019 32156
rect 58043 32100 58099 32156
rect 57963 32020 58019 32076
rect 58043 32020 58099 32076
rect 57963 31940 58019 31996
rect 58043 31940 58099 31996
rect 59206 32180 59262 32236
rect 59206 32100 59262 32156
rect 59206 32020 59262 32076
rect 59206 31940 59262 31996
rect 59364 32180 59420 32236
rect 59364 32100 59420 32156
rect 59364 32020 59420 32076
rect 59364 31940 59420 31996
rect 59672 32180 59728 32236
rect 59672 32100 59728 32156
rect 59672 32020 59728 32076
rect 59672 31940 59728 31996
rect 59818 32180 59874 32236
rect 59818 32100 59874 32156
rect 59818 32020 59874 32076
rect 59818 31940 59874 31996
rect 59954 32180 60010 32236
rect 60034 32180 60090 32236
rect 59954 32100 60010 32156
rect 60034 32100 60090 32156
rect 59954 32020 60010 32076
rect 60034 32020 60090 32076
rect 59954 31940 60010 31996
rect 60034 31940 60090 31996
rect 62326 32180 62382 32236
rect 62406 32180 62462 32236
rect 62326 32100 62382 32156
rect 62406 32100 62462 32156
rect 62326 32020 62382 32076
rect 62406 32020 62462 32076
rect 62326 31940 62382 31996
rect 62406 31940 62462 31996
rect 2044 24532 2100 24588
rect 2044 24452 2100 24508
rect 2044 24372 2100 24428
rect 2044 24292 2100 24348
rect 5540 24532 5596 24588
rect 5540 24452 5596 24508
rect 5540 24372 5596 24428
rect 5540 24292 5596 24348
rect 8430 24532 8486 24588
rect 8430 24452 8486 24508
rect 8430 24372 8486 24428
rect 8430 24292 8486 24348
rect 11320 24532 11376 24588
rect 11320 24452 11376 24508
rect 11320 24372 11376 24428
rect 11320 24292 11376 24348
rect 14210 24532 14266 24588
rect 14210 24452 14266 24508
rect 14210 24372 14266 24428
rect 14210 24292 14266 24348
rect 17100 24532 17156 24588
rect 17100 24452 17156 24508
rect 17100 24372 17156 24428
rect 17100 24292 17156 24348
rect 19990 24532 20046 24588
rect 19990 24452 20046 24508
rect 19990 24372 20046 24428
rect 19990 24292 20046 24348
rect 22880 24532 22936 24588
rect 22880 24452 22936 24508
rect 22880 24372 22936 24428
rect 22880 24292 22936 24348
rect 25770 24532 25826 24588
rect 25770 24452 25826 24508
rect 25770 24372 25826 24428
rect 25770 24292 25826 24348
rect 28660 24532 28716 24588
rect 28660 24452 28716 24508
rect 28660 24372 28716 24428
rect 28660 24292 28716 24348
rect 31550 24532 31606 24588
rect 31550 24452 31606 24508
rect 31550 24372 31606 24428
rect 31550 24292 31606 24348
rect 34440 24532 34496 24588
rect 34440 24452 34496 24508
rect 34440 24372 34496 24428
rect 34440 24292 34496 24348
rect 37330 24532 37386 24588
rect 37330 24452 37386 24508
rect 37330 24372 37386 24428
rect 37330 24292 37386 24348
rect 40220 24532 40276 24588
rect 40220 24452 40276 24508
rect 40220 24372 40276 24428
rect 40220 24292 40276 24348
rect 43110 24532 43166 24588
rect 43110 24452 43166 24508
rect 43110 24372 43166 24428
rect 43110 24292 43166 24348
rect 46000 24532 46056 24588
rect 46000 24452 46056 24508
rect 46000 24372 46056 24428
rect 46000 24292 46056 24348
rect 49008 24532 49064 24588
rect 49008 24452 49064 24508
rect 49008 24372 49064 24428
rect 49008 24292 49064 24348
rect 52237 24532 52293 24588
rect 52237 24452 52293 24508
rect 52237 24372 52293 24428
rect 52237 24292 52293 24348
rect 53638 24532 53694 24588
rect 53638 24452 53694 24508
rect 53638 24372 53694 24428
rect 53638 24292 53694 24348
rect 53806 24532 53862 24588
rect 53806 24452 53862 24508
rect 53806 24372 53862 24428
rect 53806 24292 53862 24348
rect 54550 24532 54606 24588
rect 54550 24452 54606 24508
rect 54550 24372 54606 24428
rect 54550 24292 54606 24348
rect 54940 24532 54996 24588
rect 54940 24452 54996 24508
rect 54940 24372 54996 24428
rect 54940 24292 54996 24348
rect 55656 24532 55712 24588
rect 55656 24452 55712 24508
rect 55656 24372 55712 24428
rect 55656 24292 55712 24348
rect 56234 24532 56290 24588
rect 56234 24452 56290 24508
rect 56234 24372 56290 24428
rect 56234 24292 56290 24348
rect 56679 24532 56735 24588
rect 56679 24452 56735 24508
rect 56679 24372 56735 24428
rect 56679 24292 56735 24348
rect 56983 24532 57039 24588
rect 56983 24452 57039 24508
rect 56983 24372 57039 24428
rect 56983 24292 57039 24348
rect 57825 24532 57881 24588
rect 57825 24452 57881 24508
rect 57825 24372 57881 24428
rect 57825 24292 57881 24348
rect 58465 24532 58521 24588
rect 58465 24452 58521 24508
rect 58465 24372 58521 24428
rect 58465 24292 58521 24348
rect 59048 24532 59104 24588
rect 59048 24452 59104 24508
rect 59048 24372 59104 24428
rect 59048 24292 59104 24348
rect 60326 24532 60382 24588
rect 60326 24452 60382 24508
rect 60326 24372 60382 24428
rect 60326 24292 60382 24348
rect 60484 24532 60540 24588
rect 60484 24452 60540 24508
rect 60484 24372 60540 24428
rect 60484 24292 60540 24348
rect 62528 24532 62584 24588
rect 62608 24532 62664 24588
rect 62528 24452 62584 24508
rect 62608 24452 62664 24508
rect 62528 24372 62584 24428
rect 62608 24372 62664 24428
rect 62528 24292 62584 24348
rect 62608 24292 62664 24348
rect 2184 22180 2240 22236
rect 2264 22180 2320 22236
rect 2184 22100 2240 22156
rect 2264 22100 2320 22156
rect 2184 22020 2240 22076
rect 2264 22020 2320 22076
rect 2184 21940 2240 21996
rect 2264 21940 2320 21996
rect 5393 22180 5449 22236
rect 5393 22100 5449 22156
rect 5393 22020 5449 22076
rect 5393 21940 5449 21996
rect 8283 22180 8339 22236
rect 8283 22100 8339 22156
rect 8283 22020 8339 22076
rect 8283 21940 8339 21996
rect 11173 22180 11229 22236
rect 11173 22100 11229 22156
rect 11173 22020 11229 22076
rect 11173 21940 11229 21996
rect 14063 22180 14119 22236
rect 14063 22100 14119 22156
rect 14063 22020 14119 22076
rect 14063 21940 14119 21996
rect 16953 22180 17009 22236
rect 16953 22100 17009 22156
rect 16953 22020 17009 22076
rect 16953 21940 17009 21996
rect 19843 22180 19899 22236
rect 19843 22100 19899 22156
rect 19843 22020 19899 22076
rect 19843 21940 19899 21996
rect 22733 22180 22789 22236
rect 22733 22100 22789 22156
rect 22733 22020 22789 22076
rect 22733 21940 22789 21996
rect 25623 22180 25679 22236
rect 25623 22100 25679 22156
rect 25623 22020 25679 22076
rect 25623 21940 25679 21996
rect 28513 22180 28569 22236
rect 28513 22100 28569 22156
rect 28513 22020 28569 22076
rect 28513 21940 28569 21996
rect 31403 22180 31459 22236
rect 31403 22100 31459 22156
rect 31403 22020 31459 22076
rect 31403 21940 31459 21996
rect 34293 22180 34349 22236
rect 34293 22100 34349 22156
rect 34293 22020 34349 22076
rect 34293 21940 34349 21996
rect 37183 22180 37239 22236
rect 37183 22100 37239 22156
rect 37183 22020 37239 22076
rect 37183 21940 37239 21996
rect 40073 22180 40129 22236
rect 40073 22100 40129 22156
rect 40073 22020 40129 22076
rect 40073 21940 40129 21996
rect 42963 22180 43019 22236
rect 42963 22100 43019 22156
rect 42963 22020 43019 22076
rect 42963 21940 43019 21996
rect 45853 22180 45909 22236
rect 45853 22100 45909 22156
rect 45853 22020 45909 22076
rect 45853 21940 45909 21996
rect 48800 22180 48856 22236
rect 48800 22100 48856 22156
rect 48800 22020 48856 22076
rect 48800 21940 48856 21996
rect 49662 22180 49718 22236
rect 49742 22180 49798 22236
rect 49662 22100 49718 22156
rect 49742 22100 49798 22156
rect 49662 22020 49718 22076
rect 49742 22020 49798 22076
rect 49662 21940 49718 21996
rect 49742 21940 49798 21996
rect 52956 22180 53012 22236
rect 52956 22100 53012 22156
rect 52956 22020 53012 22076
rect 52956 21940 53012 21996
rect 53114 22180 53170 22236
rect 53114 22100 53170 22156
rect 53114 22020 53170 22076
rect 53114 21940 53170 21996
rect 53470 22180 53526 22236
rect 53470 22100 53526 22156
rect 53470 22020 53526 22076
rect 53470 21940 53526 21996
rect 54788 22180 54844 22236
rect 54788 22100 54844 22156
rect 54788 22020 54844 22076
rect 54788 21940 54844 21996
rect 55381 22180 55437 22236
rect 55381 22100 55437 22156
rect 55381 22020 55437 22076
rect 55381 21940 55437 21996
rect 56527 22180 56583 22236
rect 56527 22100 56583 22156
rect 56527 22020 56583 22076
rect 56527 21940 56583 21996
rect 57963 22180 58019 22236
rect 58043 22180 58099 22236
rect 57963 22100 58019 22156
rect 58043 22100 58099 22156
rect 57963 22020 58019 22076
rect 58043 22020 58099 22076
rect 57963 21940 58019 21996
rect 58043 21940 58099 21996
rect 59206 22180 59262 22236
rect 59206 22100 59262 22156
rect 59206 22020 59262 22076
rect 59206 21940 59262 21996
rect 59364 22180 59420 22236
rect 59364 22100 59420 22156
rect 59364 22020 59420 22076
rect 59364 21940 59420 21996
rect 59672 22180 59728 22236
rect 59672 22100 59728 22156
rect 59672 22020 59728 22076
rect 59672 21940 59728 21996
rect 59818 22180 59874 22236
rect 59818 22100 59874 22156
rect 59818 22020 59874 22076
rect 59818 21940 59874 21996
rect 59954 22180 60010 22236
rect 60034 22180 60090 22236
rect 59954 22100 60010 22156
rect 60034 22100 60090 22156
rect 59954 22020 60010 22076
rect 60034 22020 60090 22076
rect 59954 21940 60010 21996
rect 60034 21940 60090 21996
rect 62326 22180 62382 22236
rect 62406 22180 62462 22236
rect 62326 22100 62382 22156
rect 62406 22100 62462 22156
rect 62326 22020 62382 22076
rect 62406 22020 62462 22076
rect 62326 21940 62382 21996
rect 62406 21940 62462 21996
rect 2044 14532 2100 14588
rect 2044 14452 2100 14508
rect 2044 14372 2100 14428
rect 2044 14292 2100 14348
rect 5540 14532 5596 14588
rect 5540 14452 5596 14508
rect 5540 14372 5596 14428
rect 5540 14292 5596 14348
rect 8430 14532 8486 14588
rect 8430 14452 8486 14508
rect 8430 14372 8486 14428
rect 8430 14292 8486 14348
rect 11320 14532 11376 14588
rect 11320 14452 11376 14508
rect 11320 14372 11376 14428
rect 11320 14292 11376 14348
rect 14210 14532 14266 14588
rect 14210 14452 14266 14508
rect 14210 14372 14266 14428
rect 14210 14292 14266 14348
rect 17100 14532 17156 14588
rect 17100 14452 17156 14508
rect 17100 14372 17156 14428
rect 17100 14292 17156 14348
rect 19990 14532 20046 14588
rect 19990 14452 20046 14508
rect 19990 14372 20046 14428
rect 19990 14292 20046 14348
rect 22880 14532 22936 14588
rect 22880 14452 22936 14508
rect 22880 14372 22936 14428
rect 22880 14292 22936 14348
rect 25770 14532 25826 14588
rect 25770 14452 25826 14508
rect 25770 14372 25826 14428
rect 25770 14292 25826 14348
rect 28660 14532 28716 14588
rect 28660 14452 28716 14508
rect 28660 14372 28716 14428
rect 28660 14292 28716 14348
rect 31550 14532 31606 14588
rect 31550 14452 31606 14508
rect 31550 14372 31606 14428
rect 31550 14292 31606 14348
rect 34440 14532 34496 14588
rect 34440 14452 34496 14508
rect 34440 14372 34496 14428
rect 34440 14292 34496 14348
rect 37330 14532 37386 14588
rect 37330 14452 37386 14508
rect 37330 14372 37386 14428
rect 37330 14292 37386 14348
rect 40220 14532 40276 14588
rect 40220 14452 40276 14508
rect 40220 14372 40276 14428
rect 40220 14292 40276 14348
rect 43110 14532 43166 14588
rect 43110 14452 43166 14508
rect 43110 14372 43166 14428
rect 43110 14292 43166 14348
rect 46000 14532 46056 14588
rect 46000 14452 46056 14508
rect 46000 14372 46056 14428
rect 46000 14292 46056 14348
rect 49008 14532 49064 14588
rect 49008 14452 49064 14508
rect 49008 14372 49064 14428
rect 49008 14292 49064 14348
rect 52237 14532 52293 14588
rect 52237 14452 52293 14508
rect 52237 14372 52293 14428
rect 52237 14292 52293 14348
rect 53638 14532 53694 14588
rect 53638 14452 53694 14508
rect 53638 14372 53694 14428
rect 53638 14292 53694 14348
rect 53806 14532 53862 14588
rect 53806 14452 53862 14508
rect 53806 14372 53862 14428
rect 53806 14292 53862 14348
rect 54550 14532 54606 14588
rect 54550 14452 54606 14508
rect 54550 14372 54606 14428
rect 54550 14292 54606 14348
rect 54940 14532 54996 14588
rect 54940 14452 54996 14508
rect 54940 14372 54996 14428
rect 54940 14292 54996 14348
rect 55656 14532 55712 14588
rect 55656 14452 55712 14508
rect 55656 14372 55712 14428
rect 55656 14292 55712 14348
rect 56234 14532 56290 14588
rect 56234 14452 56290 14508
rect 56234 14372 56290 14428
rect 56234 14292 56290 14348
rect 56679 14532 56735 14588
rect 56679 14452 56735 14508
rect 56679 14372 56735 14428
rect 56679 14292 56735 14348
rect 56983 14532 57039 14588
rect 56983 14452 57039 14508
rect 56983 14372 57039 14428
rect 56983 14292 57039 14348
rect 57825 14532 57881 14588
rect 57825 14452 57881 14508
rect 57825 14372 57881 14428
rect 57825 14292 57881 14348
rect 58465 14532 58521 14588
rect 58465 14452 58521 14508
rect 58465 14372 58521 14428
rect 58465 14292 58521 14348
rect 59048 14532 59104 14588
rect 59048 14452 59104 14508
rect 59048 14372 59104 14428
rect 59048 14292 59104 14348
rect 60326 14532 60382 14588
rect 60326 14452 60382 14508
rect 60326 14372 60382 14428
rect 60326 14292 60382 14348
rect 60484 14532 60540 14588
rect 60484 14452 60540 14508
rect 60484 14372 60540 14428
rect 60484 14292 60540 14348
rect 62528 14532 62584 14588
rect 62608 14532 62664 14588
rect 62528 14452 62584 14508
rect 62608 14452 62664 14508
rect 62528 14372 62584 14428
rect 62608 14372 62664 14428
rect 62528 14292 62584 14348
rect 62608 14292 62664 14348
rect 2184 12180 2240 12236
rect 2264 12180 2320 12236
rect 2184 12100 2240 12156
rect 2264 12100 2320 12156
rect 2184 12020 2240 12076
rect 2264 12020 2320 12076
rect 2184 11940 2240 11996
rect 2264 11940 2320 11996
rect 5393 12180 5449 12236
rect 5393 12100 5449 12156
rect 5393 12020 5449 12076
rect 5393 11940 5449 11996
rect 8283 12180 8339 12236
rect 8283 12100 8339 12156
rect 8283 12020 8339 12076
rect 8283 11940 8339 11996
rect 11173 12180 11229 12236
rect 11173 12100 11229 12156
rect 11173 12020 11229 12076
rect 11173 11940 11229 11996
rect 14063 12180 14119 12236
rect 14063 12100 14119 12156
rect 14063 12020 14119 12076
rect 14063 11940 14119 11996
rect 16953 12180 17009 12236
rect 16953 12100 17009 12156
rect 16953 12020 17009 12076
rect 16953 11940 17009 11996
rect 19843 12180 19899 12236
rect 19843 12100 19899 12156
rect 19843 12020 19899 12076
rect 19843 11940 19899 11996
rect 22733 12180 22789 12236
rect 22733 12100 22789 12156
rect 22733 12020 22789 12076
rect 22733 11940 22789 11996
rect 25623 12180 25679 12236
rect 25623 12100 25679 12156
rect 25623 12020 25679 12076
rect 25623 11940 25679 11996
rect 28513 12180 28569 12236
rect 28513 12100 28569 12156
rect 28513 12020 28569 12076
rect 28513 11940 28569 11996
rect 31403 12180 31459 12236
rect 31403 12100 31459 12156
rect 31403 12020 31459 12076
rect 31403 11940 31459 11996
rect 34293 12180 34349 12236
rect 34293 12100 34349 12156
rect 34293 12020 34349 12076
rect 34293 11940 34349 11996
rect 37183 12180 37239 12236
rect 37183 12100 37239 12156
rect 37183 12020 37239 12076
rect 37183 11940 37239 11996
rect 40073 12180 40129 12236
rect 40073 12100 40129 12156
rect 40073 12020 40129 12076
rect 40073 11940 40129 11996
rect 42963 12180 43019 12236
rect 42963 12100 43019 12156
rect 42963 12020 43019 12076
rect 42963 11940 43019 11996
rect 45853 12180 45909 12236
rect 45853 12100 45909 12156
rect 45853 12020 45909 12076
rect 45853 11940 45909 11996
rect 48800 12180 48856 12236
rect 48800 12100 48856 12156
rect 48800 12020 48856 12076
rect 48800 11940 48856 11996
rect 49662 12180 49718 12236
rect 49742 12180 49798 12236
rect 49662 12100 49718 12156
rect 49742 12100 49798 12156
rect 49662 12020 49718 12076
rect 49742 12020 49798 12076
rect 49662 11940 49718 11996
rect 49742 11940 49798 11996
rect 52956 12180 53012 12236
rect 52956 12100 53012 12156
rect 52956 12020 53012 12076
rect 52956 11940 53012 11996
rect 53114 12180 53170 12236
rect 53114 12100 53170 12156
rect 53114 12020 53170 12076
rect 53114 11940 53170 11996
rect 53470 12180 53526 12236
rect 53470 12100 53526 12156
rect 53470 12020 53526 12076
rect 53470 11940 53526 11996
rect 54788 12180 54844 12236
rect 54788 12100 54844 12156
rect 54788 12020 54844 12076
rect 54788 11940 54844 11996
rect 55381 12180 55437 12236
rect 55381 12100 55437 12156
rect 55381 12020 55437 12076
rect 55381 11940 55437 11996
rect 56527 12180 56583 12236
rect 56527 12100 56583 12156
rect 56527 12020 56583 12076
rect 56527 11940 56583 11996
rect 57963 12180 58019 12236
rect 58043 12180 58099 12236
rect 57963 12100 58019 12156
rect 58043 12100 58099 12156
rect 57963 12020 58019 12076
rect 58043 12020 58099 12076
rect 57963 11940 58019 11996
rect 58043 11940 58099 11996
rect 59206 12180 59262 12236
rect 59206 12100 59262 12156
rect 59206 12020 59262 12076
rect 59206 11940 59262 11996
rect 59364 12180 59420 12236
rect 59364 12100 59420 12156
rect 59364 12020 59420 12076
rect 59364 11940 59420 11996
rect 59672 12180 59728 12236
rect 59672 12100 59728 12156
rect 59672 12020 59728 12076
rect 59672 11940 59728 11996
rect 59818 12180 59874 12236
rect 59818 12100 59874 12156
rect 59818 12020 59874 12076
rect 59818 11940 59874 11996
rect 59954 12180 60010 12236
rect 60034 12180 60090 12236
rect 59954 12100 60010 12156
rect 60034 12100 60090 12156
rect 59954 12020 60010 12076
rect 60034 12020 60090 12076
rect 59954 11940 60010 11996
rect 60034 11940 60090 11996
rect 62326 12180 62382 12236
rect 62406 12180 62462 12236
rect 62326 12100 62382 12156
rect 62406 12100 62462 12156
rect 62326 12020 62382 12076
rect 62406 12020 62462 12076
rect 62326 11940 62382 11996
rect 62406 11940 62462 11996
rect 1864 2180 1920 2236
rect 1944 2180 2000 2236
rect 2024 2180 2080 2236
rect 2104 2180 2160 2236
rect 1864 2100 1920 2156
rect 1944 2100 2000 2156
rect 2024 2100 2080 2156
rect 2104 2100 2160 2156
rect 1864 2020 1920 2076
rect 1944 2020 2000 2076
rect 2024 2020 2080 2076
rect 2104 2020 2160 2076
rect 1864 1940 1920 1996
rect 1944 1940 2000 1996
rect 2024 1940 2080 1996
rect 2104 1940 2160 1996
rect 4216 4532 4272 4588
rect 4296 4532 4352 4588
rect 4376 4532 4432 4588
rect 4456 4532 4512 4588
rect 4216 4452 4272 4508
rect 4296 4452 4352 4508
rect 4376 4452 4432 4508
rect 4456 4452 4512 4508
rect 4216 4378 4272 4428
rect 4296 4378 4352 4428
rect 4376 4378 4432 4428
rect 4456 4378 4512 4428
rect 4216 4372 4262 4378
rect 4262 4372 4272 4378
rect 4296 4372 4326 4378
rect 4326 4372 4338 4378
rect 4338 4372 4352 4378
rect 4376 4372 4390 4378
rect 4390 4372 4402 4378
rect 4402 4372 4432 4378
rect 4456 4372 4466 4378
rect 4466 4372 4512 4378
rect 4216 4326 4262 4348
rect 4262 4326 4272 4348
rect 4296 4326 4326 4348
rect 4326 4326 4338 4348
rect 4338 4326 4352 4348
rect 4376 4326 4390 4348
rect 4390 4326 4402 4348
rect 4402 4326 4432 4348
rect 4456 4326 4466 4348
rect 4466 4326 4512 4348
rect 4216 4292 4272 4326
rect 4296 4292 4352 4326
rect 4376 4292 4432 4326
rect 4456 4292 4512 4326
rect 11864 2180 11920 2236
rect 11944 2180 12000 2236
rect 12024 2180 12080 2236
rect 12104 2180 12160 2236
rect 11864 2100 11920 2156
rect 11944 2100 12000 2156
rect 12024 2100 12080 2156
rect 12104 2100 12160 2156
rect 11864 2020 11920 2076
rect 11944 2020 12000 2076
rect 12024 2020 12080 2076
rect 12104 2020 12160 2076
rect 11864 1940 11920 1996
rect 11944 1940 12000 1996
rect 12024 1940 12080 1996
rect 12104 1940 12160 1996
rect 14216 4532 14272 4588
rect 14296 4532 14352 4588
rect 14376 4532 14432 4588
rect 14456 4532 14512 4588
rect 14216 4452 14272 4508
rect 14296 4452 14352 4508
rect 14376 4452 14432 4508
rect 14456 4452 14512 4508
rect 14216 4378 14272 4428
rect 14296 4378 14352 4428
rect 14376 4378 14432 4428
rect 14456 4378 14512 4428
rect 14216 4372 14262 4378
rect 14262 4372 14272 4378
rect 14296 4372 14326 4378
rect 14326 4372 14338 4378
rect 14338 4372 14352 4378
rect 14376 4372 14390 4378
rect 14390 4372 14402 4378
rect 14402 4372 14432 4378
rect 14456 4372 14466 4378
rect 14466 4372 14512 4378
rect 14216 4326 14262 4348
rect 14262 4326 14272 4348
rect 14296 4326 14326 4348
rect 14326 4326 14338 4348
rect 14338 4326 14352 4348
rect 14376 4326 14390 4348
rect 14390 4326 14402 4348
rect 14402 4326 14432 4348
rect 14456 4326 14466 4348
rect 14466 4326 14512 4348
rect 14216 4292 14272 4326
rect 14296 4292 14352 4326
rect 14376 4292 14432 4326
rect 14456 4292 14512 4326
rect 23018 3304 23074 3360
rect 21864 2180 21920 2236
rect 21944 2180 22000 2236
rect 22024 2180 22080 2236
rect 22104 2180 22160 2236
rect 21864 2100 21920 2156
rect 21944 2100 22000 2156
rect 22024 2100 22080 2156
rect 22104 2100 22160 2156
rect 21864 2020 21920 2076
rect 21944 2020 22000 2076
rect 22024 2020 22080 2076
rect 22104 2020 22160 2076
rect 21864 1940 21920 1996
rect 21944 1940 22000 1996
rect 22024 1940 22080 1996
rect 22104 1940 22160 1996
rect 24216 4532 24272 4588
rect 24296 4532 24352 4588
rect 24376 4532 24432 4588
rect 24456 4532 24512 4588
rect 24216 4452 24272 4508
rect 24296 4452 24352 4508
rect 24376 4452 24432 4508
rect 24456 4452 24512 4508
rect 24216 4378 24272 4428
rect 24296 4378 24352 4428
rect 24376 4378 24432 4428
rect 24456 4378 24512 4428
rect 24216 4372 24262 4378
rect 24262 4372 24272 4378
rect 24296 4372 24326 4378
rect 24326 4372 24338 4378
rect 24338 4372 24352 4378
rect 24376 4372 24390 4378
rect 24390 4372 24402 4378
rect 24402 4372 24432 4378
rect 24456 4372 24466 4378
rect 24466 4372 24512 4378
rect 24216 4326 24262 4348
rect 24262 4326 24272 4348
rect 24296 4326 24326 4348
rect 24326 4326 24338 4348
rect 24338 4326 24352 4348
rect 24376 4326 24390 4348
rect 24390 4326 24402 4348
rect 24402 4326 24432 4348
rect 24456 4326 24466 4348
rect 24466 4326 24512 4348
rect 24216 4292 24272 4326
rect 24296 4292 24352 4326
rect 24376 4292 24432 4326
rect 24456 4292 24512 4326
rect 41694 6024 41750 6080
rect 39486 5908 39542 5944
rect 39486 5888 39488 5908
rect 39488 5888 39540 5908
rect 39540 5888 39542 5908
rect 40406 5788 40408 5808
rect 40408 5788 40460 5808
rect 40460 5788 40462 5808
rect 40406 5752 40462 5788
rect 38750 5652 38752 5672
rect 38752 5652 38804 5672
rect 38804 5652 38806 5672
rect 31864 2180 31920 2236
rect 31944 2180 32000 2236
rect 32024 2180 32080 2236
rect 32104 2180 32160 2236
rect 31864 2100 31920 2156
rect 31944 2100 32000 2156
rect 32024 2100 32080 2156
rect 32104 2100 32160 2156
rect 31864 2020 31920 2076
rect 31944 2020 32000 2076
rect 32024 2020 32080 2076
rect 32104 2020 32160 2076
rect 31864 1940 31920 1996
rect 31944 1940 32000 1996
rect 32024 1940 32080 1996
rect 32104 1940 32160 1996
rect 34216 4532 34272 4588
rect 34296 4532 34352 4588
rect 34376 4532 34432 4588
rect 34456 4532 34512 4588
rect 34216 4452 34272 4508
rect 34296 4452 34352 4508
rect 34376 4452 34432 4508
rect 34456 4452 34512 4508
rect 34216 4378 34272 4428
rect 34296 4378 34352 4428
rect 34376 4378 34432 4428
rect 34456 4378 34512 4428
rect 34216 4372 34262 4378
rect 34262 4372 34272 4378
rect 34296 4372 34326 4378
rect 34326 4372 34338 4378
rect 34338 4372 34352 4378
rect 34376 4372 34390 4378
rect 34390 4372 34402 4378
rect 34402 4372 34432 4378
rect 34456 4372 34466 4378
rect 34466 4372 34512 4378
rect 34216 4326 34262 4348
rect 34262 4326 34272 4348
rect 34296 4326 34326 4348
rect 34326 4326 34338 4348
rect 34338 4326 34352 4348
rect 34376 4326 34390 4348
rect 34390 4326 34402 4348
rect 34402 4326 34432 4348
rect 34456 4326 34466 4348
rect 34466 4326 34512 4348
rect 34216 4292 34272 4326
rect 34296 4292 34352 4326
rect 34376 4292 34432 4326
rect 34456 4292 34512 4326
rect 38750 5616 38806 5652
rect 39210 5108 39212 5128
rect 39212 5108 39264 5128
rect 39264 5108 39266 5128
rect 39210 5072 39266 5108
rect 40314 3576 40370 3632
rect 40590 4800 40646 4856
rect 41326 4004 41382 4040
rect 41326 3984 41328 4004
rect 41328 3984 41380 4004
rect 41380 3984 41382 4004
rect 40866 3712 40922 3768
rect 41694 2916 41750 2952
rect 41694 2896 41696 2916
rect 41696 2896 41748 2916
rect 41748 2896 41750 2916
rect 41864 2180 41920 2236
rect 41944 2180 42000 2236
rect 42024 2180 42080 2236
rect 42104 2180 42160 2236
rect 41864 2100 41920 2156
rect 41944 2100 42000 2156
rect 42024 2100 42080 2156
rect 42104 2100 42160 2156
rect 41864 2020 41920 2076
rect 41944 2020 42000 2076
rect 42024 2020 42080 2076
rect 42104 2020 42160 2076
rect 41864 1940 41920 1996
rect 41944 1940 42000 1996
rect 42024 1940 42080 1996
rect 42104 1940 42160 1996
rect 42338 3032 42394 3088
rect 44086 5228 44142 5264
rect 44086 5208 44088 5228
rect 44088 5208 44140 5228
rect 44140 5208 44142 5228
rect 44216 4532 44272 4588
rect 44296 4532 44352 4588
rect 44376 4532 44432 4588
rect 44456 4532 44512 4588
rect 44216 4452 44272 4508
rect 44296 4452 44352 4508
rect 44376 4452 44432 4508
rect 44456 4452 44512 4508
rect 44216 4378 44272 4428
rect 44296 4378 44352 4428
rect 44376 4378 44432 4428
rect 44456 4378 44512 4428
rect 44216 4372 44262 4378
rect 44262 4372 44272 4378
rect 44296 4372 44326 4378
rect 44326 4372 44338 4378
rect 44338 4372 44352 4378
rect 44376 4372 44390 4378
rect 44390 4372 44402 4378
rect 44402 4372 44432 4378
rect 44456 4372 44466 4378
rect 44466 4372 44512 4378
rect 44216 4326 44262 4348
rect 44262 4326 44272 4348
rect 44296 4326 44326 4348
rect 44326 4326 44338 4348
rect 44338 4326 44352 4348
rect 44376 4326 44390 4348
rect 44390 4326 44402 4348
rect 44402 4326 44432 4348
rect 44456 4326 44466 4348
rect 44466 4326 44512 4348
rect 44216 4292 44272 4326
rect 44296 4292 44352 4326
rect 44376 4292 44432 4326
rect 44456 4292 44512 4326
rect 44086 3984 44142 4040
rect 42706 2896 42762 2952
rect 46202 5228 46258 5264
rect 46202 5208 46204 5228
rect 46204 5208 46256 5228
rect 46256 5208 46258 5228
rect 46662 5108 46664 5128
rect 46664 5108 46716 5128
rect 46716 5108 46718 5128
rect 46662 5072 46718 5108
rect 47582 4800 47638 4856
rect 45098 3576 45154 3632
rect 47858 3712 47914 3768
rect 47950 3032 48006 3088
rect 51262 5108 51264 5128
rect 51264 5108 51316 5128
rect 51316 5108 51318 5128
rect 51262 5072 51318 5108
rect 51864 2180 51920 2236
rect 51944 2180 52000 2236
rect 52024 2180 52080 2236
rect 52104 2180 52160 2236
rect 51864 2100 51920 2156
rect 51944 2100 52000 2156
rect 52024 2100 52080 2156
rect 52104 2100 52160 2156
rect 51864 2020 51920 2076
rect 51944 2020 52000 2076
rect 52024 2020 52080 2076
rect 52104 2020 52160 2076
rect 51864 1940 51920 1996
rect 51944 1940 52000 1996
rect 52024 1940 52080 1996
rect 52104 1940 52160 1996
rect 52826 5228 52882 5264
rect 52826 5208 52828 5228
rect 52828 5208 52880 5228
rect 52880 5208 52882 5228
rect 54850 5108 54852 5128
rect 54852 5108 54904 5128
rect 54904 5108 54906 5128
rect 54850 5072 54906 5108
rect 54216 4532 54272 4588
rect 54296 4532 54352 4588
rect 54376 4532 54432 4588
rect 54456 4532 54512 4588
rect 54216 4452 54272 4508
rect 54296 4452 54352 4508
rect 54376 4452 54432 4508
rect 54456 4452 54512 4508
rect 54216 4378 54272 4428
rect 54296 4378 54352 4428
rect 54376 4378 54432 4428
rect 54456 4378 54512 4428
rect 54216 4372 54262 4378
rect 54262 4372 54272 4378
rect 54296 4372 54326 4378
rect 54326 4372 54338 4378
rect 54338 4372 54352 4378
rect 54376 4372 54390 4378
rect 54390 4372 54402 4378
rect 54402 4372 54432 4378
rect 54456 4372 54466 4378
rect 54466 4372 54512 4378
rect 54216 4326 54262 4348
rect 54262 4326 54272 4348
rect 54296 4326 54326 4348
rect 54326 4326 54338 4348
rect 54338 4326 54352 4348
rect 54376 4326 54390 4348
rect 54390 4326 54402 4348
rect 54402 4326 54432 4348
rect 54456 4326 54466 4348
rect 54466 4326 54512 4348
rect 54216 4292 54272 4326
rect 54296 4292 54352 4326
rect 54376 4292 54432 4326
rect 54456 4292 54512 4326
rect 58530 6296 58586 6352
rect 57610 6160 57666 6216
rect 56598 5228 56654 5264
rect 56598 5208 56600 5228
rect 56600 5208 56652 5228
rect 56652 5208 56654 5228
rect 60922 6604 60924 6624
rect 60924 6604 60976 6624
rect 60976 6604 60978 6624
rect 60922 6568 60978 6604
rect 61382 6568 61438 6624
rect 61864 2180 61920 2236
rect 61944 2180 62000 2236
rect 62024 2180 62080 2236
rect 62104 2180 62160 2236
rect 61864 2100 61920 2156
rect 61944 2100 62000 2156
rect 62024 2100 62080 2156
rect 62104 2100 62160 2156
rect 61864 2020 61920 2076
rect 61944 2020 62000 2076
rect 62024 2020 62080 2076
rect 62104 2020 62160 2076
rect 61864 1940 61920 1996
rect 61944 1940 62000 1996
rect 62024 1940 62080 1996
rect 62104 1940 62160 1996
rect 62670 5888 62726 5944
rect 64142 6024 64198 6080
rect 64418 6024 64474 6080
rect 64216 4532 64272 4588
rect 64296 4532 64352 4588
rect 64376 4532 64432 4588
rect 64456 4532 64512 4588
rect 64216 4452 64272 4508
rect 64296 4452 64352 4508
rect 64376 4452 64432 4508
rect 64456 4452 64512 4508
rect 64216 4378 64272 4428
rect 64296 4378 64352 4428
rect 64376 4378 64432 4428
rect 64456 4378 64512 4428
rect 64216 4372 64262 4378
rect 64262 4372 64272 4378
rect 64296 4372 64326 4378
rect 64326 4372 64338 4378
rect 64338 4372 64352 4378
rect 64376 4372 64390 4378
rect 64390 4372 64402 4378
rect 64402 4372 64432 4378
rect 64456 4372 64466 4378
rect 64466 4372 64512 4378
rect 64216 4326 64262 4348
rect 64262 4326 64272 4348
rect 64296 4326 64326 4348
rect 64326 4326 64338 4348
rect 64338 4326 64352 4348
rect 64376 4326 64390 4348
rect 64390 4326 64402 4348
rect 64402 4326 64432 4348
rect 64456 4326 64466 4348
rect 64466 4326 64512 4348
rect 64216 4292 64272 4326
rect 64296 4292 64352 4326
rect 64376 4292 64432 4326
rect 64456 4292 64512 4326
rect 64878 7928 64934 7984
rect 65798 40976 65854 41032
rect 65430 23160 65486 23216
rect 65614 22480 65670 22536
rect 65246 7384 65302 7440
rect 65798 6332 65800 6352
rect 65800 6332 65852 6352
rect 65852 6332 65854 6352
rect 65798 6296 65854 6332
rect 65982 40160 66038 40216
rect 66626 5616 66682 5672
rect 69018 3304 69074 3360
rect 71318 6160 71374 6216
rect 71864 82180 71920 82236
rect 71944 82180 72000 82236
rect 72024 82180 72080 82236
rect 72104 82180 72160 82236
rect 71864 82118 71910 82156
rect 71910 82118 71920 82156
rect 71944 82118 71974 82156
rect 71974 82118 71986 82156
rect 71986 82118 72000 82156
rect 72024 82118 72038 82156
rect 72038 82118 72050 82156
rect 72050 82118 72080 82156
rect 72104 82118 72114 82156
rect 72114 82118 72160 82156
rect 71864 82100 71920 82118
rect 71944 82100 72000 82118
rect 72024 82100 72080 82118
rect 72104 82100 72160 82118
rect 71864 82020 71920 82076
rect 71944 82020 72000 82076
rect 72024 82020 72080 82076
rect 72104 82020 72160 82076
rect 71864 81940 71920 81996
rect 71944 81940 72000 81996
rect 72024 81940 72080 81996
rect 72104 81940 72160 81996
rect 71864 72180 71920 72236
rect 71944 72180 72000 72236
rect 72024 72180 72080 72236
rect 72104 72180 72160 72236
rect 71864 72100 71920 72156
rect 71944 72100 72000 72156
rect 72024 72100 72080 72156
rect 72104 72100 72160 72156
rect 71864 72020 71920 72076
rect 71944 72020 72000 72076
rect 72024 72020 72080 72076
rect 72104 72020 72160 72076
rect 71864 71940 71920 71996
rect 71944 71940 72000 71996
rect 72024 71940 72080 71996
rect 72104 71940 72160 71996
rect 74216 84532 74272 84588
rect 74296 84532 74352 84588
rect 74376 84532 74432 84588
rect 74456 84532 74512 84588
rect 74216 84452 74272 84508
rect 74296 84452 74352 84508
rect 74376 84452 74432 84508
rect 74456 84452 74512 84508
rect 74216 84372 74272 84428
rect 74296 84372 74352 84428
rect 74376 84372 74432 84428
rect 74456 84372 74512 84428
rect 74216 84292 74272 84348
rect 74296 84292 74352 84348
rect 74376 84292 74432 84348
rect 74456 84292 74512 84348
rect 74216 74532 74272 74588
rect 74296 74532 74352 74588
rect 74376 74532 74432 74588
rect 74456 74532 74512 74588
rect 74216 74452 74272 74508
rect 74296 74452 74352 74508
rect 74376 74452 74432 74508
rect 74456 74452 74512 74508
rect 74216 74372 74272 74428
rect 74296 74372 74352 74428
rect 74376 74372 74432 74428
rect 74456 74372 74512 74428
rect 74216 74292 74272 74348
rect 74296 74292 74352 74348
rect 74376 74292 74432 74348
rect 74456 74292 74512 74348
rect 71864 62180 71920 62236
rect 71944 62180 72000 62236
rect 72024 62180 72080 62236
rect 72104 62180 72160 62236
rect 71864 62100 71920 62156
rect 71944 62100 72000 62156
rect 72024 62100 72080 62156
rect 72104 62100 72160 62156
rect 71864 62020 71920 62076
rect 71944 62020 72000 62076
rect 72024 62020 72080 62076
rect 72104 62020 72160 62076
rect 71864 61940 71920 61996
rect 71944 61940 72000 61996
rect 72024 61940 72080 61996
rect 72104 61940 72160 61996
rect 71864 52180 71920 52236
rect 71944 52180 72000 52236
rect 72024 52180 72080 52236
rect 72104 52180 72160 52236
rect 71864 52100 71920 52156
rect 71944 52100 72000 52156
rect 72024 52100 72080 52156
rect 72104 52100 72160 52156
rect 71864 52020 71920 52076
rect 71944 52020 72000 52076
rect 72024 52020 72080 52076
rect 72104 52020 72160 52076
rect 71864 51940 71920 51996
rect 71944 51940 72000 51996
rect 72024 51940 72080 51996
rect 72104 51940 72160 51996
rect 71864 42180 71920 42236
rect 71944 42180 72000 42236
rect 72024 42180 72080 42236
rect 72104 42180 72160 42236
rect 71864 42100 71920 42156
rect 71944 42100 72000 42156
rect 72024 42100 72080 42156
rect 72104 42100 72160 42156
rect 71864 42020 71920 42076
rect 71944 42020 72000 42076
rect 72024 42020 72080 42076
rect 72104 42020 72160 42076
rect 71864 41940 71920 41996
rect 71944 41940 72000 41996
rect 72024 41940 72080 41996
rect 72104 41940 72160 41996
rect 71864 32180 71920 32236
rect 71944 32180 72000 32236
rect 72024 32180 72080 32236
rect 72104 32180 72160 32236
rect 71864 32122 71920 32156
rect 71944 32122 72000 32156
rect 72024 32122 72080 32156
rect 72104 32122 72160 32156
rect 71864 32100 71910 32122
rect 71910 32100 71920 32122
rect 71944 32100 71974 32122
rect 71974 32100 71986 32122
rect 71986 32100 72000 32122
rect 72024 32100 72038 32122
rect 72038 32100 72050 32122
rect 72050 32100 72080 32122
rect 72104 32100 72114 32122
rect 72114 32100 72160 32122
rect 71864 32070 71910 32076
rect 71910 32070 71920 32076
rect 71944 32070 71974 32076
rect 71974 32070 71986 32076
rect 71986 32070 72000 32076
rect 72024 32070 72038 32076
rect 72038 32070 72050 32076
rect 72050 32070 72080 32076
rect 72104 32070 72114 32076
rect 72114 32070 72160 32076
rect 71864 32020 71920 32070
rect 71944 32020 72000 32070
rect 72024 32020 72080 32070
rect 72104 32020 72160 32070
rect 71864 31940 71920 31996
rect 71944 31940 72000 31996
rect 72024 31940 72080 31996
rect 72104 31940 72160 31996
rect 71864 22180 71920 22236
rect 71944 22180 72000 22236
rect 72024 22180 72080 22236
rect 72104 22180 72160 22236
rect 71864 22100 71920 22156
rect 71944 22100 72000 22156
rect 72024 22100 72080 22156
rect 72104 22100 72160 22156
rect 71864 22020 71920 22076
rect 71944 22020 72000 22076
rect 72024 22020 72080 22076
rect 72104 22020 72160 22076
rect 71864 21940 71920 21996
rect 71944 21940 72000 21996
rect 72024 21940 72080 21996
rect 72104 21940 72160 21996
rect 71864 12180 71920 12236
rect 71944 12180 72000 12236
rect 72024 12180 72080 12236
rect 72104 12180 72160 12236
rect 71864 12100 71920 12156
rect 71944 12100 72000 12156
rect 72024 12100 72080 12156
rect 72104 12100 72160 12156
rect 71864 12020 71920 12076
rect 71944 12020 72000 12076
rect 72024 12020 72080 12076
rect 72104 12020 72160 12076
rect 71864 11940 71920 11996
rect 71944 11940 72000 11996
rect 72024 11940 72080 11996
rect 72104 11940 72160 11996
rect 71864 2180 71920 2236
rect 71944 2180 72000 2236
rect 72024 2180 72080 2236
rect 72104 2180 72160 2236
rect 71864 2100 71920 2156
rect 71944 2100 72000 2156
rect 72024 2100 72080 2156
rect 72104 2100 72160 2156
rect 71864 2020 71920 2076
rect 71944 2020 72000 2076
rect 72024 2020 72080 2076
rect 72104 2020 72160 2076
rect 71864 1940 71920 1996
rect 71944 1940 72000 1996
rect 72024 1940 72080 1996
rect 72104 1940 72160 1996
rect 74216 64532 74272 64588
rect 74296 64532 74352 64588
rect 74376 64532 74432 64588
rect 74456 64532 74512 64588
rect 74216 64452 74272 64508
rect 74296 64452 74352 64508
rect 74376 64452 74432 64508
rect 74456 64452 74512 64508
rect 74216 64372 74272 64428
rect 74296 64372 74352 64428
rect 74376 64372 74432 64428
rect 74456 64372 74512 64428
rect 74216 64292 74272 64348
rect 74296 64292 74352 64348
rect 74376 64292 74432 64348
rect 74456 64292 74512 64348
rect 74216 54532 74272 54588
rect 74296 54532 74352 54588
rect 74376 54532 74432 54588
rect 74456 54532 74512 54588
rect 74216 54452 74272 54508
rect 74296 54452 74352 54508
rect 74376 54452 74432 54508
rect 74456 54452 74512 54508
rect 74216 54426 74272 54428
rect 74296 54426 74352 54428
rect 74376 54426 74432 54428
rect 74456 54426 74512 54428
rect 74216 54374 74262 54426
rect 74262 54374 74272 54426
rect 74296 54374 74326 54426
rect 74326 54374 74338 54426
rect 74338 54374 74352 54426
rect 74376 54374 74390 54426
rect 74390 54374 74402 54426
rect 74402 54374 74432 54426
rect 74456 54374 74466 54426
rect 74466 54374 74512 54426
rect 74216 54372 74272 54374
rect 74296 54372 74352 54374
rect 74376 54372 74432 54374
rect 74456 54372 74512 54374
rect 74216 54292 74272 54348
rect 74296 54292 74352 54348
rect 74376 54292 74432 54348
rect 74456 54292 74512 54348
rect 74216 44582 74262 44588
rect 74262 44582 74272 44588
rect 74296 44582 74326 44588
rect 74326 44582 74338 44588
rect 74338 44582 74352 44588
rect 74376 44582 74390 44588
rect 74390 44582 74402 44588
rect 74402 44582 74432 44588
rect 74456 44582 74466 44588
rect 74466 44582 74512 44588
rect 74216 44532 74272 44582
rect 74296 44532 74352 44582
rect 74376 44532 74432 44582
rect 74456 44532 74512 44582
rect 74216 44452 74272 44508
rect 74296 44452 74352 44508
rect 74376 44452 74432 44508
rect 74456 44452 74512 44508
rect 74216 44372 74272 44428
rect 74296 44372 74352 44428
rect 74376 44372 74432 44428
rect 74456 44372 74512 44428
rect 74216 44292 74272 44348
rect 74296 44292 74352 44348
rect 74376 44292 74432 44348
rect 74456 44292 74512 44348
rect 74216 34532 74272 34588
rect 74296 34532 74352 34588
rect 74376 34532 74432 34588
rect 74456 34532 74512 34588
rect 74216 34452 74272 34508
rect 74296 34452 74352 34508
rect 74376 34452 74432 34508
rect 74456 34452 74512 34508
rect 74216 34372 74272 34428
rect 74296 34372 74352 34428
rect 74376 34372 74432 34428
rect 74456 34372 74512 34428
rect 74216 34292 74272 34348
rect 74296 34292 74352 34348
rect 74376 34292 74432 34348
rect 74456 34292 74512 34348
rect 74216 24532 74272 24588
rect 74296 24532 74352 24588
rect 74376 24532 74432 24588
rect 74456 24532 74512 24588
rect 74216 24452 74272 24508
rect 74296 24452 74352 24508
rect 74376 24452 74432 24508
rect 74456 24452 74512 24508
rect 74216 24372 74272 24428
rect 74296 24372 74352 24428
rect 74376 24372 74432 24428
rect 74456 24372 74512 24428
rect 74216 24292 74272 24348
rect 74296 24292 74352 24348
rect 74376 24292 74432 24348
rect 74456 24292 74512 24348
rect 74216 14532 74272 14588
rect 74296 14532 74352 14588
rect 74376 14532 74432 14588
rect 74456 14532 74512 14588
rect 74216 14452 74272 14508
rect 74296 14452 74352 14508
rect 74376 14452 74432 14508
rect 74456 14452 74512 14508
rect 74216 14372 74272 14428
rect 74296 14372 74352 14428
rect 74376 14372 74432 14428
rect 74456 14372 74512 14428
rect 74216 14292 74272 14348
rect 74296 14292 74352 14348
rect 74376 14292 74432 14348
rect 74456 14292 74512 14348
rect 74216 4532 74272 4588
rect 74296 4532 74352 4588
rect 74376 4532 74432 4588
rect 74456 4532 74512 4588
rect 74216 4452 74272 4508
rect 74296 4452 74352 4508
rect 74376 4452 74432 4508
rect 74456 4452 74512 4508
rect 74216 4378 74272 4428
rect 74296 4378 74352 4428
rect 74376 4378 74432 4428
rect 74456 4378 74512 4428
rect 74216 4372 74262 4378
rect 74262 4372 74272 4378
rect 74296 4372 74326 4378
rect 74326 4372 74338 4378
rect 74338 4372 74352 4378
rect 74376 4372 74390 4378
rect 74390 4372 74402 4378
rect 74402 4372 74432 4378
rect 74456 4372 74466 4378
rect 74466 4372 74512 4378
rect 74216 4326 74262 4348
rect 74262 4326 74272 4348
rect 74296 4326 74326 4348
rect 74326 4326 74338 4348
rect 74338 4326 74352 4348
rect 74376 4326 74390 4348
rect 74390 4326 74402 4348
rect 74402 4326 74432 4348
rect 74456 4326 74466 4348
rect 74466 4326 74512 4348
rect 74216 4292 74272 4326
rect 74296 4292 74352 4326
rect 74376 4292 74432 4326
rect 74456 4292 74512 4326
<< metal3 >>
rect 964 84588 75028 84616
rect 964 84532 2044 84588
rect 2100 84532 5540 84588
rect 5596 84532 8430 84588
rect 8486 84532 11320 84588
rect 11376 84532 14210 84588
rect 14266 84532 17100 84588
rect 17156 84532 19990 84588
rect 20046 84532 22880 84588
rect 22936 84532 25770 84588
rect 25826 84532 28660 84588
rect 28716 84532 31550 84588
rect 31606 84532 34440 84588
rect 34496 84532 37330 84588
rect 37386 84532 40220 84588
rect 40276 84532 43110 84588
rect 43166 84532 46000 84588
rect 46056 84532 49008 84588
rect 49064 84532 52237 84588
rect 52293 84532 53638 84588
rect 53694 84532 53806 84588
rect 53862 84532 54550 84588
rect 54606 84532 54940 84588
rect 54996 84532 55656 84588
rect 55712 84532 56234 84588
rect 56290 84532 56679 84588
rect 56735 84532 56983 84588
rect 57039 84532 57825 84588
rect 57881 84532 58465 84588
rect 58521 84532 59048 84588
rect 59104 84532 60326 84588
rect 60382 84532 60484 84588
rect 60540 84532 62528 84588
rect 62584 84532 62608 84588
rect 62664 84532 74216 84588
rect 74272 84532 74296 84588
rect 74352 84532 74376 84588
rect 74432 84532 74456 84588
rect 74512 84532 75028 84588
rect 964 84508 75028 84532
rect 964 84452 2044 84508
rect 2100 84452 5540 84508
rect 5596 84452 8430 84508
rect 8486 84452 11320 84508
rect 11376 84452 14210 84508
rect 14266 84452 17100 84508
rect 17156 84452 19990 84508
rect 20046 84452 22880 84508
rect 22936 84452 25770 84508
rect 25826 84452 28660 84508
rect 28716 84452 31550 84508
rect 31606 84452 34440 84508
rect 34496 84452 37330 84508
rect 37386 84452 40220 84508
rect 40276 84452 43110 84508
rect 43166 84452 46000 84508
rect 46056 84452 49008 84508
rect 49064 84452 52237 84508
rect 52293 84452 53638 84508
rect 53694 84452 53806 84508
rect 53862 84452 54550 84508
rect 54606 84452 54940 84508
rect 54996 84452 55656 84508
rect 55712 84452 56234 84508
rect 56290 84452 56679 84508
rect 56735 84452 56983 84508
rect 57039 84452 57825 84508
rect 57881 84452 58465 84508
rect 58521 84452 59048 84508
rect 59104 84452 60326 84508
rect 60382 84452 60484 84508
rect 60540 84452 62528 84508
rect 62584 84452 62608 84508
rect 62664 84452 74216 84508
rect 74272 84452 74296 84508
rect 74352 84452 74376 84508
rect 74432 84452 74456 84508
rect 74512 84452 75028 84508
rect 964 84428 75028 84452
rect 964 84372 2044 84428
rect 2100 84372 5540 84428
rect 5596 84372 8430 84428
rect 8486 84372 11320 84428
rect 11376 84372 14210 84428
rect 14266 84372 17100 84428
rect 17156 84372 19990 84428
rect 20046 84372 22880 84428
rect 22936 84372 25770 84428
rect 25826 84372 28660 84428
rect 28716 84372 31550 84428
rect 31606 84372 34440 84428
rect 34496 84372 37330 84428
rect 37386 84372 40220 84428
rect 40276 84372 43110 84428
rect 43166 84372 46000 84428
rect 46056 84372 49008 84428
rect 49064 84372 52237 84428
rect 52293 84372 53638 84428
rect 53694 84372 53806 84428
rect 53862 84372 54550 84428
rect 54606 84372 54940 84428
rect 54996 84372 55656 84428
rect 55712 84372 56234 84428
rect 56290 84372 56679 84428
rect 56735 84372 56983 84428
rect 57039 84372 57825 84428
rect 57881 84372 58465 84428
rect 58521 84372 59048 84428
rect 59104 84372 60326 84428
rect 60382 84372 60484 84428
rect 60540 84372 62528 84428
rect 62584 84372 62608 84428
rect 62664 84372 74216 84428
rect 74272 84372 74296 84428
rect 74352 84372 74376 84428
rect 74432 84372 74456 84428
rect 74512 84372 75028 84428
rect 964 84348 75028 84372
rect 964 84292 2044 84348
rect 2100 84292 5540 84348
rect 5596 84292 8430 84348
rect 8486 84292 11320 84348
rect 11376 84292 14210 84348
rect 14266 84292 17100 84348
rect 17156 84292 19990 84348
rect 20046 84292 22880 84348
rect 22936 84292 25770 84348
rect 25826 84292 28660 84348
rect 28716 84292 31550 84348
rect 31606 84292 34440 84348
rect 34496 84292 37330 84348
rect 37386 84292 40220 84348
rect 40276 84292 43110 84348
rect 43166 84292 46000 84348
rect 46056 84292 49008 84348
rect 49064 84292 52237 84348
rect 52293 84292 53638 84348
rect 53694 84292 53806 84348
rect 53862 84292 54550 84348
rect 54606 84292 54940 84348
rect 54996 84292 55656 84348
rect 55712 84292 56234 84348
rect 56290 84292 56679 84348
rect 56735 84292 56983 84348
rect 57039 84292 57825 84348
rect 57881 84292 58465 84348
rect 58521 84292 59048 84348
rect 59104 84292 60326 84348
rect 60382 84292 60484 84348
rect 60540 84292 62528 84348
rect 62584 84292 62608 84348
rect 62664 84292 74216 84348
rect 74272 84292 74296 84348
rect 74352 84292 74376 84348
rect 74432 84292 74456 84348
rect 74512 84292 75028 84348
rect 964 84264 75028 84292
rect 964 82236 75028 82264
rect 964 82180 2184 82236
rect 2240 82180 2264 82236
rect 2320 82180 5393 82236
rect 5449 82180 8283 82236
rect 8339 82180 11173 82236
rect 11229 82180 14063 82236
rect 14119 82180 16953 82236
rect 17009 82180 19843 82236
rect 19899 82180 22733 82236
rect 22789 82180 25623 82236
rect 25679 82180 28513 82236
rect 28569 82180 31403 82236
rect 31459 82180 34293 82236
rect 34349 82180 37183 82236
rect 37239 82180 40073 82236
rect 40129 82180 42963 82236
rect 43019 82180 45853 82236
rect 45909 82180 48800 82236
rect 48856 82180 49662 82236
rect 49718 82180 49742 82236
rect 49798 82180 52956 82236
rect 53012 82180 53114 82236
rect 53170 82180 53470 82236
rect 53526 82180 54788 82236
rect 54844 82180 55381 82236
rect 55437 82180 56527 82236
rect 56583 82180 57963 82236
rect 58019 82180 58043 82236
rect 58099 82180 59206 82236
rect 59262 82180 59364 82236
rect 59420 82180 59672 82236
rect 59728 82180 59818 82236
rect 59874 82180 59954 82236
rect 60010 82180 60034 82236
rect 60090 82180 62326 82236
rect 62382 82180 62406 82236
rect 62462 82180 71864 82236
rect 71920 82180 71944 82236
rect 72000 82180 72024 82236
rect 72080 82180 72104 82236
rect 72160 82180 75028 82236
rect 964 82156 75028 82180
rect 964 82100 2184 82156
rect 2240 82100 2264 82156
rect 2320 82100 5393 82156
rect 5449 82100 8283 82156
rect 8339 82100 11173 82156
rect 11229 82100 14063 82156
rect 14119 82100 16953 82156
rect 17009 82100 19843 82156
rect 19899 82100 22733 82156
rect 22789 82100 25623 82156
rect 25679 82100 28513 82156
rect 28569 82100 31403 82156
rect 31459 82100 34293 82156
rect 34349 82100 37183 82156
rect 37239 82100 40073 82156
rect 40129 82100 42963 82156
rect 43019 82100 45853 82156
rect 45909 82100 48800 82156
rect 48856 82100 49662 82156
rect 49718 82100 49742 82156
rect 49798 82100 52956 82156
rect 53012 82100 53114 82156
rect 53170 82100 53470 82156
rect 53526 82100 54788 82156
rect 54844 82100 55381 82156
rect 55437 82100 56527 82156
rect 56583 82100 57963 82156
rect 58019 82100 58043 82156
rect 58099 82100 59206 82156
rect 59262 82100 59364 82156
rect 59420 82100 59672 82156
rect 59728 82100 59818 82156
rect 59874 82100 59954 82156
rect 60010 82100 60034 82156
rect 60090 82100 62326 82156
rect 62382 82100 62406 82156
rect 62462 82100 71864 82156
rect 71920 82100 71944 82156
rect 72000 82100 72024 82156
rect 72080 82100 72104 82156
rect 72160 82100 75028 82156
rect 964 82076 75028 82100
rect 964 82020 2184 82076
rect 2240 82020 2264 82076
rect 2320 82020 5393 82076
rect 5449 82020 8283 82076
rect 8339 82020 11173 82076
rect 11229 82020 14063 82076
rect 14119 82020 16953 82076
rect 17009 82020 19843 82076
rect 19899 82020 22733 82076
rect 22789 82020 25623 82076
rect 25679 82020 28513 82076
rect 28569 82020 31403 82076
rect 31459 82020 34293 82076
rect 34349 82020 37183 82076
rect 37239 82020 40073 82076
rect 40129 82020 42963 82076
rect 43019 82020 45853 82076
rect 45909 82020 48800 82076
rect 48856 82020 49662 82076
rect 49718 82020 49742 82076
rect 49798 82020 52956 82076
rect 53012 82020 53114 82076
rect 53170 82020 53470 82076
rect 53526 82020 54788 82076
rect 54844 82020 55381 82076
rect 55437 82020 56527 82076
rect 56583 82020 57963 82076
rect 58019 82020 58043 82076
rect 58099 82020 59206 82076
rect 59262 82020 59364 82076
rect 59420 82020 59672 82076
rect 59728 82020 59818 82076
rect 59874 82020 59954 82076
rect 60010 82020 60034 82076
rect 60090 82020 62326 82076
rect 62382 82020 62406 82076
rect 62462 82020 71864 82076
rect 71920 82020 71944 82076
rect 72000 82020 72024 82076
rect 72080 82020 72104 82076
rect 72160 82020 75028 82076
rect 964 81996 75028 82020
rect 964 81940 2184 81996
rect 2240 81940 2264 81996
rect 2320 81940 5393 81996
rect 5449 81940 8283 81996
rect 8339 81940 11173 81996
rect 11229 81940 14063 81996
rect 14119 81940 16953 81996
rect 17009 81940 19843 81996
rect 19899 81940 22733 81996
rect 22789 81940 25623 81996
rect 25679 81940 28513 81996
rect 28569 81940 31403 81996
rect 31459 81940 34293 81996
rect 34349 81940 37183 81996
rect 37239 81940 40073 81996
rect 40129 81940 42963 81996
rect 43019 81940 45853 81996
rect 45909 81940 48800 81996
rect 48856 81940 49662 81996
rect 49718 81940 49742 81996
rect 49798 81940 52956 81996
rect 53012 81940 53114 81996
rect 53170 81940 53470 81996
rect 53526 81940 54788 81996
rect 54844 81940 55381 81996
rect 55437 81940 56527 81996
rect 56583 81940 57963 81996
rect 58019 81940 58043 81996
rect 58099 81940 59206 81996
rect 59262 81940 59364 81996
rect 59420 81940 59672 81996
rect 59728 81940 59818 81996
rect 59874 81940 59954 81996
rect 60010 81940 60034 81996
rect 60090 81940 62326 81996
rect 62382 81940 62406 81996
rect 62462 81940 71864 81996
rect 71920 81940 71944 81996
rect 72000 81940 72024 81996
rect 72080 81940 72104 81996
rect 72160 81940 75028 81996
rect 964 81912 75028 81940
rect 964 74588 75028 74616
rect 964 74532 2044 74588
rect 2100 74532 5540 74588
rect 5596 74532 8430 74588
rect 8486 74532 11320 74588
rect 11376 74532 14210 74588
rect 14266 74532 17100 74588
rect 17156 74532 19990 74588
rect 20046 74532 22880 74588
rect 22936 74532 25770 74588
rect 25826 74532 28660 74588
rect 28716 74532 31550 74588
rect 31606 74532 34440 74588
rect 34496 74532 37330 74588
rect 37386 74532 40220 74588
rect 40276 74532 43110 74588
rect 43166 74532 46000 74588
rect 46056 74532 49008 74588
rect 49064 74532 52237 74588
rect 52293 74532 53638 74588
rect 53694 74532 53806 74588
rect 53862 74532 54550 74588
rect 54606 74532 54940 74588
rect 54996 74532 55656 74588
rect 55712 74532 56234 74588
rect 56290 74532 56679 74588
rect 56735 74532 56983 74588
rect 57039 74532 57825 74588
rect 57881 74532 58465 74588
rect 58521 74532 59048 74588
rect 59104 74532 60326 74588
rect 60382 74532 60484 74588
rect 60540 74532 62528 74588
rect 62584 74532 62608 74588
rect 62664 74532 74216 74588
rect 74272 74532 74296 74588
rect 74352 74532 74376 74588
rect 74432 74532 74456 74588
rect 74512 74532 75028 74588
rect 964 74508 75028 74532
rect 964 74452 2044 74508
rect 2100 74452 5540 74508
rect 5596 74452 8430 74508
rect 8486 74452 11320 74508
rect 11376 74452 14210 74508
rect 14266 74452 17100 74508
rect 17156 74452 19990 74508
rect 20046 74452 22880 74508
rect 22936 74452 25770 74508
rect 25826 74452 28660 74508
rect 28716 74452 31550 74508
rect 31606 74452 34440 74508
rect 34496 74452 37330 74508
rect 37386 74452 40220 74508
rect 40276 74452 43110 74508
rect 43166 74452 46000 74508
rect 46056 74452 49008 74508
rect 49064 74452 52237 74508
rect 52293 74452 53638 74508
rect 53694 74452 53806 74508
rect 53862 74452 54550 74508
rect 54606 74452 54940 74508
rect 54996 74452 55656 74508
rect 55712 74452 56234 74508
rect 56290 74452 56679 74508
rect 56735 74452 56983 74508
rect 57039 74452 57825 74508
rect 57881 74452 58465 74508
rect 58521 74452 59048 74508
rect 59104 74452 60326 74508
rect 60382 74452 60484 74508
rect 60540 74452 62528 74508
rect 62584 74452 62608 74508
rect 62664 74452 74216 74508
rect 74272 74452 74296 74508
rect 74352 74452 74376 74508
rect 74432 74452 74456 74508
rect 74512 74452 75028 74508
rect 964 74428 75028 74452
rect 964 74372 2044 74428
rect 2100 74372 5540 74428
rect 5596 74372 8430 74428
rect 8486 74372 11320 74428
rect 11376 74372 14210 74428
rect 14266 74372 17100 74428
rect 17156 74372 19990 74428
rect 20046 74372 22880 74428
rect 22936 74372 25770 74428
rect 25826 74372 28660 74428
rect 28716 74372 31550 74428
rect 31606 74372 34440 74428
rect 34496 74372 37330 74428
rect 37386 74372 40220 74428
rect 40276 74372 43110 74428
rect 43166 74372 46000 74428
rect 46056 74372 49008 74428
rect 49064 74372 52237 74428
rect 52293 74372 53638 74428
rect 53694 74372 53806 74428
rect 53862 74372 54550 74428
rect 54606 74372 54940 74428
rect 54996 74372 55656 74428
rect 55712 74372 56234 74428
rect 56290 74372 56679 74428
rect 56735 74372 56983 74428
rect 57039 74372 57825 74428
rect 57881 74372 58465 74428
rect 58521 74372 59048 74428
rect 59104 74372 60326 74428
rect 60382 74372 60484 74428
rect 60540 74372 62528 74428
rect 62584 74372 62608 74428
rect 62664 74372 74216 74428
rect 74272 74372 74296 74428
rect 74352 74372 74376 74428
rect 74432 74372 74456 74428
rect 74512 74372 75028 74428
rect 964 74348 75028 74372
rect 964 74292 2044 74348
rect 2100 74292 5540 74348
rect 5596 74292 8430 74348
rect 8486 74292 11320 74348
rect 11376 74292 14210 74348
rect 14266 74292 17100 74348
rect 17156 74292 19990 74348
rect 20046 74292 22880 74348
rect 22936 74292 25770 74348
rect 25826 74292 28660 74348
rect 28716 74292 31550 74348
rect 31606 74292 34440 74348
rect 34496 74292 37330 74348
rect 37386 74292 40220 74348
rect 40276 74292 43110 74348
rect 43166 74292 46000 74348
rect 46056 74292 49008 74348
rect 49064 74292 52237 74348
rect 52293 74292 53638 74348
rect 53694 74292 53806 74348
rect 53862 74292 54550 74348
rect 54606 74292 54940 74348
rect 54996 74292 55656 74348
rect 55712 74292 56234 74348
rect 56290 74292 56679 74348
rect 56735 74292 56983 74348
rect 57039 74292 57825 74348
rect 57881 74292 58465 74348
rect 58521 74292 59048 74348
rect 59104 74292 60326 74348
rect 60382 74292 60484 74348
rect 60540 74292 62528 74348
rect 62584 74292 62608 74348
rect 62664 74292 74216 74348
rect 74272 74292 74296 74348
rect 74352 74292 74376 74348
rect 74432 74292 74456 74348
rect 74512 74292 75028 74348
rect 964 74264 75028 74292
rect 964 72236 75028 72264
rect 964 72180 2184 72236
rect 2240 72180 2264 72236
rect 2320 72180 5393 72236
rect 5449 72180 8283 72236
rect 8339 72180 11173 72236
rect 11229 72180 14063 72236
rect 14119 72180 16953 72236
rect 17009 72180 19843 72236
rect 19899 72180 22733 72236
rect 22789 72180 25623 72236
rect 25679 72180 28513 72236
rect 28569 72180 31403 72236
rect 31459 72180 34293 72236
rect 34349 72180 37183 72236
rect 37239 72180 40073 72236
rect 40129 72180 42963 72236
rect 43019 72180 45853 72236
rect 45909 72180 48800 72236
rect 48856 72180 49662 72236
rect 49718 72180 49742 72236
rect 49798 72180 52956 72236
rect 53012 72180 53114 72236
rect 53170 72180 53470 72236
rect 53526 72180 54788 72236
rect 54844 72180 55381 72236
rect 55437 72180 56527 72236
rect 56583 72180 57963 72236
rect 58019 72180 58043 72236
rect 58099 72180 59206 72236
rect 59262 72180 59364 72236
rect 59420 72180 59672 72236
rect 59728 72180 59818 72236
rect 59874 72180 59954 72236
rect 60010 72180 60034 72236
rect 60090 72180 62326 72236
rect 62382 72180 62406 72236
rect 62462 72180 71864 72236
rect 71920 72180 71944 72236
rect 72000 72180 72024 72236
rect 72080 72180 72104 72236
rect 72160 72180 75028 72236
rect 964 72156 75028 72180
rect 964 72100 2184 72156
rect 2240 72100 2264 72156
rect 2320 72100 5393 72156
rect 5449 72100 8283 72156
rect 8339 72100 11173 72156
rect 11229 72100 14063 72156
rect 14119 72100 16953 72156
rect 17009 72100 19843 72156
rect 19899 72100 22733 72156
rect 22789 72100 25623 72156
rect 25679 72100 28513 72156
rect 28569 72100 31403 72156
rect 31459 72100 34293 72156
rect 34349 72100 37183 72156
rect 37239 72100 40073 72156
rect 40129 72100 42963 72156
rect 43019 72100 45853 72156
rect 45909 72100 48800 72156
rect 48856 72100 49662 72156
rect 49718 72100 49742 72156
rect 49798 72100 52956 72156
rect 53012 72100 53114 72156
rect 53170 72100 53470 72156
rect 53526 72100 54788 72156
rect 54844 72100 55381 72156
rect 55437 72100 56527 72156
rect 56583 72100 57963 72156
rect 58019 72100 58043 72156
rect 58099 72100 59206 72156
rect 59262 72100 59364 72156
rect 59420 72100 59672 72156
rect 59728 72100 59818 72156
rect 59874 72100 59954 72156
rect 60010 72100 60034 72156
rect 60090 72100 62326 72156
rect 62382 72100 62406 72156
rect 62462 72100 71864 72156
rect 71920 72100 71944 72156
rect 72000 72100 72024 72156
rect 72080 72100 72104 72156
rect 72160 72100 75028 72156
rect 964 72076 75028 72100
rect 964 72020 2184 72076
rect 2240 72020 2264 72076
rect 2320 72020 5393 72076
rect 5449 72020 8283 72076
rect 8339 72020 11173 72076
rect 11229 72020 14063 72076
rect 14119 72020 16953 72076
rect 17009 72020 19843 72076
rect 19899 72020 22733 72076
rect 22789 72020 25623 72076
rect 25679 72020 28513 72076
rect 28569 72020 31403 72076
rect 31459 72020 34293 72076
rect 34349 72020 37183 72076
rect 37239 72020 40073 72076
rect 40129 72020 42963 72076
rect 43019 72020 45853 72076
rect 45909 72020 48800 72076
rect 48856 72020 49662 72076
rect 49718 72020 49742 72076
rect 49798 72020 52956 72076
rect 53012 72020 53114 72076
rect 53170 72020 53470 72076
rect 53526 72020 54788 72076
rect 54844 72020 55381 72076
rect 55437 72020 56527 72076
rect 56583 72020 57963 72076
rect 58019 72020 58043 72076
rect 58099 72020 59206 72076
rect 59262 72020 59364 72076
rect 59420 72020 59672 72076
rect 59728 72020 59818 72076
rect 59874 72020 59954 72076
rect 60010 72020 60034 72076
rect 60090 72020 62326 72076
rect 62382 72020 62406 72076
rect 62462 72020 71864 72076
rect 71920 72020 71944 72076
rect 72000 72020 72024 72076
rect 72080 72020 72104 72076
rect 72160 72020 75028 72076
rect 964 71996 75028 72020
rect 964 71940 2184 71996
rect 2240 71940 2264 71996
rect 2320 71940 5393 71996
rect 5449 71940 8283 71996
rect 8339 71940 11173 71996
rect 11229 71940 14063 71996
rect 14119 71940 16953 71996
rect 17009 71940 19843 71996
rect 19899 71940 22733 71996
rect 22789 71940 25623 71996
rect 25679 71940 28513 71996
rect 28569 71940 31403 71996
rect 31459 71940 34293 71996
rect 34349 71940 37183 71996
rect 37239 71940 40073 71996
rect 40129 71940 42963 71996
rect 43019 71940 45853 71996
rect 45909 71940 48800 71996
rect 48856 71940 49662 71996
rect 49718 71940 49742 71996
rect 49798 71940 52956 71996
rect 53012 71940 53114 71996
rect 53170 71940 53470 71996
rect 53526 71940 54788 71996
rect 54844 71940 55381 71996
rect 55437 71940 56527 71996
rect 56583 71940 57963 71996
rect 58019 71940 58043 71996
rect 58099 71940 59206 71996
rect 59262 71940 59364 71996
rect 59420 71940 59672 71996
rect 59728 71940 59818 71996
rect 59874 71940 59954 71996
rect 60010 71940 60034 71996
rect 60090 71940 62326 71996
rect 62382 71940 62406 71996
rect 62462 71940 71864 71996
rect 71920 71940 71944 71996
rect 72000 71940 72024 71996
rect 72080 71940 72104 71996
rect 72160 71940 75028 71996
rect 964 71912 75028 71940
rect 964 64588 75028 64616
rect 964 64532 2044 64588
rect 2100 64532 5540 64588
rect 5596 64532 8430 64588
rect 8486 64532 11320 64588
rect 11376 64532 14210 64588
rect 14266 64532 17100 64588
rect 17156 64532 19990 64588
rect 20046 64532 22880 64588
rect 22936 64532 25770 64588
rect 25826 64532 28660 64588
rect 28716 64532 31550 64588
rect 31606 64532 34440 64588
rect 34496 64532 37330 64588
rect 37386 64532 40220 64588
rect 40276 64532 43110 64588
rect 43166 64532 46000 64588
rect 46056 64532 49008 64588
rect 49064 64532 52237 64588
rect 52293 64532 53638 64588
rect 53694 64532 53806 64588
rect 53862 64532 54550 64588
rect 54606 64532 54940 64588
rect 54996 64532 55656 64588
rect 55712 64532 56234 64588
rect 56290 64532 56679 64588
rect 56735 64532 56983 64588
rect 57039 64532 57825 64588
rect 57881 64532 58465 64588
rect 58521 64532 59048 64588
rect 59104 64532 60326 64588
rect 60382 64532 60484 64588
rect 60540 64532 62528 64588
rect 62584 64532 62608 64588
rect 62664 64532 74216 64588
rect 74272 64532 74296 64588
rect 74352 64532 74376 64588
rect 74432 64532 74456 64588
rect 74512 64532 75028 64588
rect 964 64508 75028 64532
rect 964 64452 2044 64508
rect 2100 64452 5540 64508
rect 5596 64452 8430 64508
rect 8486 64452 11320 64508
rect 11376 64452 14210 64508
rect 14266 64452 17100 64508
rect 17156 64452 19990 64508
rect 20046 64452 22880 64508
rect 22936 64452 25770 64508
rect 25826 64452 28660 64508
rect 28716 64452 31550 64508
rect 31606 64452 34440 64508
rect 34496 64452 37330 64508
rect 37386 64452 40220 64508
rect 40276 64452 43110 64508
rect 43166 64452 46000 64508
rect 46056 64452 49008 64508
rect 49064 64452 52237 64508
rect 52293 64452 53638 64508
rect 53694 64452 53806 64508
rect 53862 64452 54550 64508
rect 54606 64452 54940 64508
rect 54996 64452 55656 64508
rect 55712 64452 56234 64508
rect 56290 64452 56679 64508
rect 56735 64452 56983 64508
rect 57039 64452 57825 64508
rect 57881 64452 58465 64508
rect 58521 64452 59048 64508
rect 59104 64452 60326 64508
rect 60382 64452 60484 64508
rect 60540 64452 62528 64508
rect 62584 64452 62608 64508
rect 62664 64452 74216 64508
rect 74272 64452 74296 64508
rect 74352 64452 74376 64508
rect 74432 64452 74456 64508
rect 74512 64452 75028 64508
rect 964 64428 75028 64452
rect 964 64372 2044 64428
rect 2100 64372 5540 64428
rect 5596 64372 8430 64428
rect 8486 64372 11320 64428
rect 11376 64372 14210 64428
rect 14266 64372 17100 64428
rect 17156 64372 19990 64428
rect 20046 64372 22880 64428
rect 22936 64372 25770 64428
rect 25826 64372 28660 64428
rect 28716 64372 31550 64428
rect 31606 64372 34440 64428
rect 34496 64372 37330 64428
rect 37386 64372 40220 64428
rect 40276 64372 43110 64428
rect 43166 64372 46000 64428
rect 46056 64372 49008 64428
rect 49064 64372 52237 64428
rect 52293 64372 53638 64428
rect 53694 64372 53806 64428
rect 53862 64372 54550 64428
rect 54606 64372 54940 64428
rect 54996 64372 55656 64428
rect 55712 64372 56234 64428
rect 56290 64372 56679 64428
rect 56735 64372 56983 64428
rect 57039 64372 57825 64428
rect 57881 64372 58465 64428
rect 58521 64372 59048 64428
rect 59104 64372 60326 64428
rect 60382 64372 60484 64428
rect 60540 64372 62528 64428
rect 62584 64372 62608 64428
rect 62664 64372 74216 64428
rect 74272 64372 74296 64428
rect 74352 64372 74376 64428
rect 74432 64372 74456 64428
rect 74512 64372 75028 64428
rect 964 64348 75028 64372
rect 964 64292 2044 64348
rect 2100 64292 5540 64348
rect 5596 64292 8430 64348
rect 8486 64292 11320 64348
rect 11376 64292 14210 64348
rect 14266 64292 17100 64348
rect 17156 64292 19990 64348
rect 20046 64292 22880 64348
rect 22936 64292 25770 64348
rect 25826 64292 28660 64348
rect 28716 64292 31550 64348
rect 31606 64292 34440 64348
rect 34496 64292 37330 64348
rect 37386 64292 40220 64348
rect 40276 64292 43110 64348
rect 43166 64292 46000 64348
rect 46056 64292 49008 64348
rect 49064 64292 52237 64348
rect 52293 64292 53638 64348
rect 53694 64292 53806 64348
rect 53862 64292 54550 64348
rect 54606 64292 54940 64348
rect 54996 64292 55656 64348
rect 55712 64292 56234 64348
rect 56290 64292 56679 64348
rect 56735 64292 56983 64348
rect 57039 64292 57825 64348
rect 57881 64292 58465 64348
rect 58521 64292 59048 64348
rect 59104 64292 60326 64348
rect 60382 64292 60484 64348
rect 60540 64292 62528 64348
rect 62584 64292 62608 64348
rect 62664 64292 74216 64348
rect 74272 64292 74296 64348
rect 74352 64292 74376 64348
rect 74432 64292 74456 64348
rect 74512 64292 75028 64348
rect 964 64264 75028 64292
rect 964 62236 75028 62264
rect 964 62180 2184 62236
rect 2240 62180 2264 62236
rect 2320 62180 5393 62236
rect 5449 62180 8283 62236
rect 8339 62180 11173 62236
rect 11229 62180 14063 62236
rect 14119 62180 16953 62236
rect 17009 62180 19843 62236
rect 19899 62180 22733 62236
rect 22789 62180 25623 62236
rect 25679 62180 28513 62236
rect 28569 62180 31403 62236
rect 31459 62180 34293 62236
rect 34349 62180 37183 62236
rect 37239 62180 40073 62236
rect 40129 62180 42963 62236
rect 43019 62180 45853 62236
rect 45909 62180 48800 62236
rect 48856 62180 49662 62236
rect 49718 62180 49742 62236
rect 49798 62180 52956 62236
rect 53012 62180 53114 62236
rect 53170 62180 53470 62236
rect 53526 62180 54788 62236
rect 54844 62180 55381 62236
rect 55437 62180 56527 62236
rect 56583 62180 57963 62236
rect 58019 62180 58043 62236
rect 58099 62180 59206 62236
rect 59262 62180 59364 62236
rect 59420 62180 59672 62236
rect 59728 62180 59818 62236
rect 59874 62180 59954 62236
rect 60010 62180 60034 62236
rect 60090 62180 62326 62236
rect 62382 62180 62406 62236
rect 62462 62180 71864 62236
rect 71920 62180 71944 62236
rect 72000 62180 72024 62236
rect 72080 62180 72104 62236
rect 72160 62180 75028 62236
rect 964 62156 75028 62180
rect 964 62100 2184 62156
rect 2240 62100 2264 62156
rect 2320 62100 5393 62156
rect 5449 62100 8283 62156
rect 8339 62100 11173 62156
rect 11229 62100 14063 62156
rect 14119 62100 16953 62156
rect 17009 62100 19843 62156
rect 19899 62100 22733 62156
rect 22789 62100 25623 62156
rect 25679 62100 28513 62156
rect 28569 62100 31403 62156
rect 31459 62100 34293 62156
rect 34349 62100 37183 62156
rect 37239 62100 40073 62156
rect 40129 62100 42963 62156
rect 43019 62100 45853 62156
rect 45909 62100 48800 62156
rect 48856 62100 49662 62156
rect 49718 62100 49742 62156
rect 49798 62100 52956 62156
rect 53012 62100 53114 62156
rect 53170 62100 53470 62156
rect 53526 62100 54788 62156
rect 54844 62100 55381 62156
rect 55437 62100 56527 62156
rect 56583 62100 57963 62156
rect 58019 62100 58043 62156
rect 58099 62100 59206 62156
rect 59262 62100 59364 62156
rect 59420 62100 59672 62156
rect 59728 62100 59818 62156
rect 59874 62100 59954 62156
rect 60010 62100 60034 62156
rect 60090 62100 62326 62156
rect 62382 62100 62406 62156
rect 62462 62100 71864 62156
rect 71920 62100 71944 62156
rect 72000 62100 72024 62156
rect 72080 62100 72104 62156
rect 72160 62100 75028 62156
rect 964 62076 75028 62100
rect 964 62020 2184 62076
rect 2240 62020 2264 62076
rect 2320 62020 5393 62076
rect 5449 62020 8283 62076
rect 8339 62020 11173 62076
rect 11229 62020 14063 62076
rect 14119 62020 16953 62076
rect 17009 62020 19843 62076
rect 19899 62020 22733 62076
rect 22789 62020 25623 62076
rect 25679 62020 28513 62076
rect 28569 62020 31403 62076
rect 31459 62020 34293 62076
rect 34349 62020 37183 62076
rect 37239 62020 40073 62076
rect 40129 62020 42963 62076
rect 43019 62020 45853 62076
rect 45909 62020 48800 62076
rect 48856 62020 49662 62076
rect 49718 62020 49742 62076
rect 49798 62020 52956 62076
rect 53012 62020 53114 62076
rect 53170 62020 53470 62076
rect 53526 62020 54788 62076
rect 54844 62020 55381 62076
rect 55437 62020 56527 62076
rect 56583 62020 57963 62076
rect 58019 62020 58043 62076
rect 58099 62020 59206 62076
rect 59262 62020 59364 62076
rect 59420 62020 59672 62076
rect 59728 62020 59818 62076
rect 59874 62020 59954 62076
rect 60010 62020 60034 62076
rect 60090 62020 62326 62076
rect 62382 62020 62406 62076
rect 62462 62020 71864 62076
rect 71920 62020 71944 62076
rect 72000 62020 72024 62076
rect 72080 62020 72104 62076
rect 72160 62020 75028 62076
rect 964 61996 75028 62020
rect 964 61940 2184 61996
rect 2240 61940 2264 61996
rect 2320 61940 5393 61996
rect 5449 61940 8283 61996
rect 8339 61940 11173 61996
rect 11229 61940 14063 61996
rect 14119 61940 16953 61996
rect 17009 61940 19843 61996
rect 19899 61940 22733 61996
rect 22789 61940 25623 61996
rect 25679 61940 28513 61996
rect 28569 61940 31403 61996
rect 31459 61940 34293 61996
rect 34349 61940 37183 61996
rect 37239 61940 40073 61996
rect 40129 61940 42963 61996
rect 43019 61940 45853 61996
rect 45909 61940 48800 61996
rect 48856 61940 49662 61996
rect 49718 61940 49742 61996
rect 49798 61940 52956 61996
rect 53012 61940 53114 61996
rect 53170 61940 53470 61996
rect 53526 61940 54788 61996
rect 54844 61940 55381 61996
rect 55437 61940 56527 61996
rect 56583 61940 57963 61996
rect 58019 61940 58043 61996
rect 58099 61940 59206 61996
rect 59262 61940 59364 61996
rect 59420 61940 59672 61996
rect 59728 61940 59818 61996
rect 59874 61940 59954 61996
rect 60010 61940 60034 61996
rect 60090 61940 62326 61996
rect 62382 61940 62406 61996
rect 62462 61940 71864 61996
rect 71920 61940 71944 61996
rect 72000 61940 72024 61996
rect 72080 61940 72104 61996
rect 72160 61940 75028 61996
rect 964 61912 75028 61940
rect 964 54588 75028 54616
rect 964 54532 2044 54588
rect 2100 54532 5540 54588
rect 5596 54532 8430 54588
rect 8486 54532 11320 54588
rect 11376 54532 14210 54588
rect 14266 54532 17100 54588
rect 17156 54532 19990 54588
rect 20046 54532 22880 54588
rect 22936 54532 25770 54588
rect 25826 54532 28660 54588
rect 28716 54532 31550 54588
rect 31606 54532 34440 54588
rect 34496 54532 37330 54588
rect 37386 54532 40220 54588
rect 40276 54532 43110 54588
rect 43166 54532 46000 54588
rect 46056 54532 49008 54588
rect 49064 54532 52237 54588
rect 52293 54532 53638 54588
rect 53694 54532 53806 54588
rect 53862 54532 54550 54588
rect 54606 54532 54940 54588
rect 54996 54532 55656 54588
rect 55712 54532 56234 54588
rect 56290 54532 56679 54588
rect 56735 54532 56983 54588
rect 57039 54532 57825 54588
rect 57881 54532 58465 54588
rect 58521 54532 59048 54588
rect 59104 54532 60326 54588
rect 60382 54532 60484 54588
rect 60540 54532 62528 54588
rect 62584 54532 62608 54588
rect 62664 54532 74216 54588
rect 74272 54532 74296 54588
rect 74352 54532 74376 54588
rect 74432 54532 74456 54588
rect 74512 54532 75028 54588
rect 964 54508 75028 54532
rect 964 54452 2044 54508
rect 2100 54452 5540 54508
rect 5596 54452 8430 54508
rect 8486 54452 11320 54508
rect 11376 54452 14210 54508
rect 14266 54452 17100 54508
rect 17156 54452 19990 54508
rect 20046 54452 22880 54508
rect 22936 54452 25770 54508
rect 25826 54452 28660 54508
rect 28716 54452 31550 54508
rect 31606 54452 34440 54508
rect 34496 54452 37330 54508
rect 37386 54452 40220 54508
rect 40276 54452 43110 54508
rect 43166 54452 46000 54508
rect 46056 54452 49008 54508
rect 49064 54452 52237 54508
rect 52293 54452 53638 54508
rect 53694 54452 53806 54508
rect 53862 54452 54550 54508
rect 54606 54452 54940 54508
rect 54996 54452 55656 54508
rect 55712 54452 56234 54508
rect 56290 54452 56679 54508
rect 56735 54452 56983 54508
rect 57039 54452 57825 54508
rect 57881 54452 58465 54508
rect 58521 54452 59048 54508
rect 59104 54452 60326 54508
rect 60382 54452 60484 54508
rect 60540 54452 62528 54508
rect 62584 54452 62608 54508
rect 62664 54452 74216 54508
rect 74272 54452 74296 54508
rect 74352 54452 74376 54508
rect 74432 54452 74456 54508
rect 74512 54452 75028 54508
rect 964 54428 75028 54452
rect 964 54372 2044 54428
rect 2100 54372 5540 54428
rect 5596 54372 8430 54428
rect 8486 54372 11320 54428
rect 11376 54372 14210 54428
rect 14266 54372 17100 54428
rect 17156 54372 19990 54428
rect 20046 54372 22880 54428
rect 22936 54372 25770 54428
rect 25826 54372 28660 54428
rect 28716 54372 31550 54428
rect 31606 54372 34440 54428
rect 34496 54372 37330 54428
rect 37386 54372 40220 54428
rect 40276 54372 43110 54428
rect 43166 54372 46000 54428
rect 46056 54372 49008 54428
rect 49064 54372 52237 54428
rect 52293 54372 53638 54428
rect 53694 54372 53806 54428
rect 53862 54372 54550 54428
rect 54606 54372 54940 54428
rect 54996 54372 55656 54428
rect 55712 54372 56234 54428
rect 56290 54372 56679 54428
rect 56735 54372 56983 54428
rect 57039 54372 57825 54428
rect 57881 54372 58465 54428
rect 58521 54372 59048 54428
rect 59104 54372 60326 54428
rect 60382 54372 60484 54428
rect 60540 54372 62528 54428
rect 62584 54372 62608 54428
rect 62664 54372 74216 54428
rect 74272 54372 74296 54428
rect 74352 54372 74376 54428
rect 74432 54372 74456 54428
rect 74512 54372 75028 54428
rect 964 54348 75028 54372
rect 964 54292 2044 54348
rect 2100 54292 5540 54348
rect 5596 54292 8430 54348
rect 8486 54292 11320 54348
rect 11376 54292 14210 54348
rect 14266 54292 17100 54348
rect 17156 54292 19990 54348
rect 20046 54292 22880 54348
rect 22936 54292 25770 54348
rect 25826 54292 28660 54348
rect 28716 54292 31550 54348
rect 31606 54292 34440 54348
rect 34496 54292 37330 54348
rect 37386 54292 40220 54348
rect 40276 54292 43110 54348
rect 43166 54292 46000 54348
rect 46056 54292 49008 54348
rect 49064 54292 52237 54348
rect 52293 54292 53638 54348
rect 53694 54292 53806 54348
rect 53862 54292 54550 54348
rect 54606 54292 54940 54348
rect 54996 54292 55656 54348
rect 55712 54292 56234 54348
rect 56290 54292 56679 54348
rect 56735 54292 56983 54348
rect 57039 54292 57825 54348
rect 57881 54292 58465 54348
rect 58521 54292 59048 54348
rect 59104 54292 60326 54348
rect 60382 54292 60484 54348
rect 60540 54292 62528 54348
rect 62584 54292 62608 54348
rect 62664 54292 74216 54348
rect 74272 54292 74296 54348
rect 74352 54292 74376 54348
rect 74432 54292 74456 54348
rect 74512 54292 75028 54348
rect 964 54264 75028 54292
rect 964 52236 75028 52264
rect 964 52180 2184 52236
rect 2240 52180 2264 52236
rect 2320 52180 5393 52236
rect 5449 52180 8283 52236
rect 8339 52180 11173 52236
rect 11229 52180 14063 52236
rect 14119 52180 16953 52236
rect 17009 52180 19843 52236
rect 19899 52180 22733 52236
rect 22789 52180 25623 52236
rect 25679 52180 28513 52236
rect 28569 52180 31403 52236
rect 31459 52180 34293 52236
rect 34349 52180 37183 52236
rect 37239 52180 40073 52236
rect 40129 52180 42963 52236
rect 43019 52180 45853 52236
rect 45909 52180 48800 52236
rect 48856 52180 49662 52236
rect 49718 52180 49742 52236
rect 49798 52180 52956 52236
rect 53012 52180 53114 52236
rect 53170 52180 53470 52236
rect 53526 52180 54788 52236
rect 54844 52180 55381 52236
rect 55437 52180 56527 52236
rect 56583 52180 57963 52236
rect 58019 52180 58043 52236
rect 58099 52180 59206 52236
rect 59262 52180 59364 52236
rect 59420 52180 59672 52236
rect 59728 52180 59818 52236
rect 59874 52180 59954 52236
rect 60010 52180 60034 52236
rect 60090 52180 62326 52236
rect 62382 52180 62406 52236
rect 62462 52180 71864 52236
rect 71920 52180 71944 52236
rect 72000 52180 72024 52236
rect 72080 52180 72104 52236
rect 72160 52180 75028 52236
rect 964 52156 75028 52180
rect 964 52100 2184 52156
rect 2240 52100 2264 52156
rect 2320 52100 5393 52156
rect 5449 52100 8283 52156
rect 8339 52100 11173 52156
rect 11229 52100 14063 52156
rect 14119 52100 16953 52156
rect 17009 52100 19843 52156
rect 19899 52100 22733 52156
rect 22789 52100 25623 52156
rect 25679 52100 28513 52156
rect 28569 52100 31403 52156
rect 31459 52100 34293 52156
rect 34349 52100 37183 52156
rect 37239 52100 40073 52156
rect 40129 52100 42963 52156
rect 43019 52100 45853 52156
rect 45909 52100 48800 52156
rect 48856 52100 49662 52156
rect 49718 52100 49742 52156
rect 49798 52100 52956 52156
rect 53012 52100 53114 52156
rect 53170 52100 53470 52156
rect 53526 52100 54788 52156
rect 54844 52100 55381 52156
rect 55437 52100 56527 52156
rect 56583 52100 57963 52156
rect 58019 52100 58043 52156
rect 58099 52100 59206 52156
rect 59262 52100 59364 52156
rect 59420 52100 59672 52156
rect 59728 52100 59818 52156
rect 59874 52100 59954 52156
rect 60010 52100 60034 52156
rect 60090 52100 62326 52156
rect 62382 52100 62406 52156
rect 62462 52100 71864 52156
rect 71920 52100 71944 52156
rect 72000 52100 72024 52156
rect 72080 52100 72104 52156
rect 72160 52100 75028 52156
rect 964 52076 75028 52100
rect 964 52020 2184 52076
rect 2240 52020 2264 52076
rect 2320 52020 5393 52076
rect 5449 52020 8283 52076
rect 8339 52020 11173 52076
rect 11229 52020 14063 52076
rect 14119 52020 16953 52076
rect 17009 52020 19843 52076
rect 19899 52020 22733 52076
rect 22789 52020 25623 52076
rect 25679 52020 28513 52076
rect 28569 52020 31403 52076
rect 31459 52020 34293 52076
rect 34349 52020 37183 52076
rect 37239 52020 40073 52076
rect 40129 52020 42963 52076
rect 43019 52020 45853 52076
rect 45909 52020 48800 52076
rect 48856 52020 49662 52076
rect 49718 52020 49742 52076
rect 49798 52020 52956 52076
rect 53012 52020 53114 52076
rect 53170 52020 53470 52076
rect 53526 52020 54788 52076
rect 54844 52020 55381 52076
rect 55437 52020 56527 52076
rect 56583 52020 57963 52076
rect 58019 52020 58043 52076
rect 58099 52020 59206 52076
rect 59262 52020 59364 52076
rect 59420 52020 59672 52076
rect 59728 52020 59818 52076
rect 59874 52020 59954 52076
rect 60010 52020 60034 52076
rect 60090 52020 62326 52076
rect 62382 52020 62406 52076
rect 62462 52020 71864 52076
rect 71920 52020 71944 52076
rect 72000 52020 72024 52076
rect 72080 52020 72104 52076
rect 72160 52020 75028 52076
rect 964 51996 75028 52020
rect 964 51940 2184 51996
rect 2240 51940 2264 51996
rect 2320 51940 5393 51996
rect 5449 51940 8283 51996
rect 8339 51940 11173 51996
rect 11229 51940 14063 51996
rect 14119 51940 16953 51996
rect 17009 51940 19843 51996
rect 19899 51940 22733 51996
rect 22789 51940 25623 51996
rect 25679 51940 28513 51996
rect 28569 51940 31403 51996
rect 31459 51940 34293 51996
rect 34349 51940 37183 51996
rect 37239 51940 40073 51996
rect 40129 51940 42963 51996
rect 43019 51940 45853 51996
rect 45909 51940 48800 51996
rect 48856 51940 49662 51996
rect 49718 51940 49742 51996
rect 49798 51940 52956 51996
rect 53012 51940 53114 51996
rect 53170 51940 53470 51996
rect 53526 51940 54788 51996
rect 54844 51940 55381 51996
rect 55437 51940 56527 51996
rect 56583 51940 57963 51996
rect 58019 51940 58043 51996
rect 58099 51940 59206 51996
rect 59262 51940 59364 51996
rect 59420 51940 59672 51996
rect 59728 51940 59818 51996
rect 59874 51940 59954 51996
rect 60010 51940 60034 51996
rect 60090 51940 62326 51996
rect 62382 51940 62406 51996
rect 62462 51940 71864 51996
rect 71920 51940 71944 51996
rect 72000 51940 72024 51996
rect 72080 51940 72104 51996
rect 72160 51940 75028 51996
rect 964 51912 75028 51940
rect 964 44588 75028 44616
rect 964 44532 2044 44588
rect 2100 44532 5540 44588
rect 5596 44532 8430 44588
rect 8486 44532 11320 44588
rect 11376 44532 14210 44588
rect 14266 44532 17100 44588
rect 17156 44532 19990 44588
rect 20046 44532 22880 44588
rect 22936 44532 25770 44588
rect 25826 44532 28660 44588
rect 28716 44532 31550 44588
rect 31606 44532 34440 44588
rect 34496 44532 37330 44588
rect 37386 44532 40220 44588
rect 40276 44532 43110 44588
rect 43166 44532 46000 44588
rect 46056 44532 52237 44588
rect 52293 44532 53638 44588
rect 53694 44532 54550 44588
rect 54606 44532 54940 44588
rect 54996 44532 55656 44588
rect 55712 44532 56234 44588
rect 56290 44532 56679 44588
rect 56735 44532 56983 44588
rect 57039 44532 57825 44588
rect 57881 44532 58349 44588
rect 58405 44532 59048 44588
rect 59104 44532 60326 44588
rect 60382 44532 60484 44588
rect 60540 44532 62528 44588
rect 62584 44532 62608 44588
rect 62664 44532 74216 44588
rect 74272 44532 74296 44588
rect 74352 44532 74376 44588
rect 74432 44532 74456 44588
rect 74512 44532 75028 44588
rect 964 44508 75028 44532
rect 964 44452 2044 44508
rect 2100 44452 5540 44508
rect 5596 44452 8430 44508
rect 8486 44452 11320 44508
rect 11376 44452 14210 44508
rect 14266 44452 17100 44508
rect 17156 44452 19990 44508
rect 20046 44452 22880 44508
rect 22936 44452 25770 44508
rect 25826 44452 28660 44508
rect 28716 44452 31550 44508
rect 31606 44452 34440 44508
rect 34496 44452 37330 44508
rect 37386 44452 40220 44508
rect 40276 44452 43110 44508
rect 43166 44452 46000 44508
rect 46056 44452 52237 44508
rect 52293 44452 53638 44508
rect 53694 44452 54550 44508
rect 54606 44452 54940 44508
rect 54996 44452 55656 44508
rect 55712 44452 56234 44508
rect 56290 44452 56679 44508
rect 56735 44452 56983 44508
rect 57039 44452 57825 44508
rect 57881 44452 58349 44508
rect 58405 44452 59048 44508
rect 59104 44452 60326 44508
rect 60382 44452 60484 44508
rect 60540 44452 62528 44508
rect 62584 44452 62608 44508
rect 62664 44452 74216 44508
rect 74272 44452 74296 44508
rect 74352 44452 74376 44508
rect 74432 44452 74456 44508
rect 74512 44452 75028 44508
rect 964 44428 75028 44452
rect 964 44372 2044 44428
rect 2100 44372 5540 44428
rect 5596 44372 8430 44428
rect 8486 44372 11320 44428
rect 11376 44372 14210 44428
rect 14266 44372 17100 44428
rect 17156 44372 19990 44428
rect 20046 44372 22880 44428
rect 22936 44372 25770 44428
rect 25826 44372 28660 44428
rect 28716 44372 31550 44428
rect 31606 44372 34440 44428
rect 34496 44372 37330 44428
rect 37386 44372 40220 44428
rect 40276 44372 43110 44428
rect 43166 44372 46000 44428
rect 46056 44372 52237 44428
rect 52293 44372 53638 44428
rect 53694 44372 54550 44428
rect 54606 44372 54940 44428
rect 54996 44372 55656 44428
rect 55712 44372 56234 44428
rect 56290 44372 56679 44428
rect 56735 44372 56983 44428
rect 57039 44372 57825 44428
rect 57881 44372 58349 44428
rect 58405 44372 59048 44428
rect 59104 44372 60326 44428
rect 60382 44372 60484 44428
rect 60540 44372 62528 44428
rect 62584 44372 62608 44428
rect 62664 44372 74216 44428
rect 74272 44372 74296 44428
rect 74352 44372 74376 44428
rect 74432 44372 74456 44428
rect 74512 44372 75028 44428
rect 964 44348 75028 44372
rect 964 44292 2044 44348
rect 2100 44292 5540 44348
rect 5596 44292 8430 44348
rect 8486 44292 11320 44348
rect 11376 44292 14210 44348
rect 14266 44292 17100 44348
rect 17156 44292 19990 44348
rect 20046 44292 22880 44348
rect 22936 44292 25770 44348
rect 25826 44292 28660 44348
rect 28716 44292 31550 44348
rect 31606 44292 34440 44348
rect 34496 44292 37330 44348
rect 37386 44292 40220 44348
rect 40276 44292 43110 44348
rect 43166 44292 46000 44348
rect 46056 44292 52237 44348
rect 52293 44292 53638 44348
rect 53694 44292 54550 44348
rect 54606 44292 54940 44348
rect 54996 44292 55656 44348
rect 55712 44292 56234 44348
rect 56290 44292 56679 44348
rect 56735 44292 56983 44348
rect 57039 44292 57825 44348
rect 57881 44292 58349 44348
rect 58405 44292 59048 44348
rect 59104 44292 60326 44348
rect 60382 44292 60484 44348
rect 60540 44292 62528 44348
rect 62584 44292 62608 44348
rect 62664 44292 74216 44348
rect 74272 44292 74296 44348
rect 74352 44292 74376 44348
rect 74432 44292 74456 44348
rect 74512 44292 75028 44348
rect 964 44264 75028 44292
rect 964 42236 75028 42264
rect 964 42180 2184 42236
rect 2240 42180 2264 42236
rect 2320 42180 5393 42236
rect 5449 42180 8283 42236
rect 8339 42180 11173 42236
rect 11229 42180 14063 42236
rect 14119 42180 16953 42236
rect 17009 42180 19843 42236
rect 19899 42180 22733 42236
rect 22789 42180 25623 42236
rect 25679 42180 28513 42236
rect 28569 42180 31403 42236
rect 31459 42180 34293 42236
rect 34349 42180 37183 42236
rect 37239 42180 40073 42236
rect 40129 42180 42963 42236
rect 43019 42180 45853 42236
rect 45909 42180 48800 42236
rect 48856 42180 49662 42236
rect 49718 42180 49742 42236
rect 49798 42180 52956 42236
rect 53012 42180 53114 42236
rect 53170 42180 53470 42236
rect 53526 42180 54788 42236
rect 54844 42180 55381 42236
rect 55437 42180 56527 42236
rect 56583 42180 57963 42236
rect 58019 42180 58043 42236
rect 58099 42180 59206 42236
rect 59262 42180 59364 42236
rect 59420 42180 59672 42236
rect 59728 42180 59818 42236
rect 59874 42180 59954 42236
rect 60010 42180 60034 42236
rect 60090 42180 62326 42236
rect 62382 42180 62406 42236
rect 62462 42180 71864 42236
rect 71920 42180 71944 42236
rect 72000 42180 72024 42236
rect 72080 42180 72104 42236
rect 72160 42180 75028 42236
rect 964 42156 75028 42180
rect 964 42100 2184 42156
rect 2240 42100 2264 42156
rect 2320 42100 5393 42156
rect 5449 42100 8283 42156
rect 8339 42100 11173 42156
rect 11229 42100 14063 42156
rect 14119 42100 16953 42156
rect 17009 42100 19843 42156
rect 19899 42100 22733 42156
rect 22789 42100 25623 42156
rect 25679 42100 28513 42156
rect 28569 42100 31403 42156
rect 31459 42100 34293 42156
rect 34349 42100 37183 42156
rect 37239 42100 40073 42156
rect 40129 42100 42963 42156
rect 43019 42100 45853 42156
rect 45909 42100 48800 42156
rect 48856 42100 49662 42156
rect 49718 42100 49742 42156
rect 49798 42100 52956 42156
rect 53012 42100 53114 42156
rect 53170 42100 53470 42156
rect 53526 42100 54788 42156
rect 54844 42100 55381 42156
rect 55437 42100 56527 42156
rect 56583 42100 57963 42156
rect 58019 42100 58043 42156
rect 58099 42100 59206 42156
rect 59262 42100 59364 42156
rect 59420 42100 59672 42156
rect 59728 42100 59818 42156
rect 59874 42100 59954 42156
rect 60010 42100 60034 42156
rect 60090 42100 62326 42156
rect 62382 42100 62406 42156
rect 62462 42100 71864 42156
rect 71920 42100 71944 42156
rect 72000 42100 72024 42156
rect 72080 42100 72104 42156
rect 72160 42100 75028 42156
rect 964 42076 75028 42100
rect 964 42020 2184 42076
rect 2240 42020 2264 42076
rect 2320 42020 5393 42076
rect 5449 42020 8283 42076
rect 8339 42020 11173 42076
rect 11229 42020 14063 42076
rect 14119 42020 16953 42076
rect 17009 42020 19843 42076
rect 19899 42020 22733 42076
rect 22789 42020 25623 42076
rect 25679 42020 28513 42076
rect 28569 42020 31403 42076
rect 31459 42020 34293 42076
rect 34349 42020 37183 42076
rect 37239 42020 40073 42076
rect 40129 42020 42963 42076
rect 43019 42020 45853 42076
rect 45909 42020 48800 42076
rect 48856 42020 49662 42076
rect 49718 42020 49742 42076
rect 49798 42020 52956 42076
rect 53012 42020 53114 42076
rect 53170 42020 53470 42076
rect 53526 42020 54788 42076
rect 54844 42020 55381 42076
rect 55437 42020 56527 42076
rect 56583 42020 57963 42076
rect 58019 42020 58043 42076
rect 58099 42020 59206 42076
rect 59262 42020 59364 42076
rect 59420 42020 59672 42076
rect 59728 42020 59818 42076
rect 59874 42020 59954 42076
rect 60010 42020 60034 42076
rect 60090 42020 62326 42076
rect 62382 42020 62406 42076
rect 62462 42020 71864 42076
rect 71920 42020 71944 42076
rect 72000 42020 72024 42076
rect 72080 42020 72104 42076
rect 72160 42020 75028 42076
rect 964 41996 75028 42020
rect 964 41940 2184 41996
rect 2240 41940 2264 41996
rect 2320 41940 5393 41996
rect 5449 41940 8283 41996
rect 8339 41940 11173 41996
rect 11229 41940 14063 41996
rect 14119 41940 16953 41996
rect 17009 41940 19843 41996
rect 19899 41940 22733 41996
rect 22789 41940 25623 41996
rect 25679 41940 28513 41996
rect 28569 41940 31403 41996
rect 31459 41940 34293 41996
rect 34349 41940 37183 41996
rect 37239 41940 40073 41996
rect 40129 41940 42963 41996
rect 43019 41940 45853 41996
rect 45909 41940 48800 41996
rect 48856 41940 49662 41996
rect 49718 41940 49742 41996
rect 49798 41940 52956 41996
rect 53012 41940 53114 41996
rect 53170 41940 53470 41996
rect 53526 41940 54788 41996
rect 54844 41940 55381 41996
rect 55437 41940 56527 41996
rect 56583 41940 57963 41996
rect 58019 41940 58043 41996
rect 58099 41940 59206 41996
rect 59262 41940 59364 41996
rect 59420 41940 59672 41996
rect 59728 41940 59818 41996
rect 59874 41940 59954 41996
rect 60010 41940 60034 41996
rect 60090 41940 62326 41996
rect 62382 41940 62406 41996
rect 62462 41940 71864 41996
rect 71920 41940 71944 41996
rect 72000 41940 72024 41996
rect 72080 41940 72104 41996
rect 72160 41940 75028 41996
rect 964 41912 75028 41940
rect 65793 41034 65859 41037
rect 65793 41032 65994 41034
rect 65793 40976 65798 41032
rect 65854 40976 65994 41032
rect 65793 40974 65994 40976
rect 65793 40971 65859 40974
rect 65934 40221 65994 40974
rect 65934 40216 66043 40221
rect 65934 40160 65982 40216
rect 66038 40160 66043 40216
rect 65934 40158 66043 40160
rect 65977 40155 66043 40158
rect 964 34588 75028 34616
rect 964 34532 2044 34588
rect 2100 34532 5540 34588
rect 5596 34532 8430 34588
rect 8486 34532 11320 34588
rect 11376 34532 14210 34588
rect 14266 34532 17100 34588
rect 17156 34532 19990 34588
rect 20046 34532 22880 34588
rect 22936 34532 25770 34588
rect 25826 34532 28660 34588
rect 28716 34532 31550 34588
rect 31606 34532 34440 34588
rect 34496 34532 37330 34588
rect 37386 34532 40220 34588
rect 40276 34532 43110 34588
rect 43166 34532 46000 34588
rect 46056 34532 49008 34588
rect 49064 34532 52237 34588
rect 52293 34532 53638 34588
rect 53694 34532 53806 34588
rect 53862 34532 54550 34588
rect 54606 34532 54940 34588
rect 54996 34532 55656 34588
rect 55712 34532 56234 34588
rect 56290 34532 56679 34588
rect 56735 34532 56983 34588
rect 57039 34532 57825 34588
rect 57881 34532 58465 34588
rect 58521 34532 59048 34588
rect 59104 34532 60326 34588
rect 60382 34532 60484 34588
rect 60540 34532 62528 34588
rect 62584 34532 62608 34588
rect 62664 34532 74216 34588
rect 74272 34532 74296 34588
rect 74352 34532 74376 34588
rect 74432 34532 74456 34588
rect 74512 34532 75028 34588
rect 964 34508 75028 34532
rect 964 34452 2044 34508
rect 2100 34452 5540 34508
rect 5596 34452 8430 34508
rect 8486 34452 11320 34508
rect 11376 34452 14210 34508
rect 14266 34452 17100 34508
rect 17156 34452 19990 34508
rect 20046 34452 22880 34508
rect 22936 34452 25770 34508
rect 25826 34452 28660 34508
rect 28716 34452 31550 34508
rect 31606 34452 34440 34508
rect 34496 34452 37330 34508
rect 37386 34452 40220 34508
rect 40276 34452 43110 34508
rect 43166 34452 46000 34508
rect 46056 34452 49008 34508
rect 49064 34452 52237 34508
rect 52293 34452 53638 34508
rect 53694 34452 53806 34508
rect 53862 34452 54550 34508
rect 54606 34452 54940 34508
rect 54996 34452 55656 34508
rect 55712 34452 56234 34508
rect 56290 34452 56679 34508
rect 56735 34452 56983 34508
rect 57039 34452 57825 34508
rect 57881 34452 58465 34508
rect 58521 34452 59048 34508
rect 59104 34452 60326 34508
rect 60382 34452 60484 34508
rect 60540 34452 62528 34508
rect 62584 34452 62608 34508
rect 62664 34452 74216 34508
rect 74272 34452 74296 34508
rect 74352 34452 74376 34508
rect 74432 34452 74456 34508
rect 74512 34452 75028 34508
rect 964 34428 75028 34452
rect 964 34372 2044 34428
rect 2100 34372 5540 34428
rect 5596 34372 8430 34428
rect 8486 34372 11320 34428
rect 11376 34372 14210 34428
rect 14266 34372 17100 34428
rect 17156 34372 19990 34428
rect 20046 34372 22880 34428
rect 22936 34372 25770 34428
rect 25826 34372 28660 34428
rect 28716 34372 31550 34428
rect 31606 34372 34440 34428
rect 34496 34372 37330 34428
rect 37386 34372 40220 34428
rect 40276 34372 43110 34428
rect 43166 34372 46000 34428
rect 46056 34372 49008 34428
rect 49064 34372 52237 34428
rect 52293 34372 53638 34428
rect 53694 34372 53806 34428
rect 53862 34372 54550 34428
rect 54606 34372 54940 34428
rect 54996 34372 55656 34428
rect 55712 34372 56234 34428
rect 56290 34372 56679 34428
rect 56735 34372 56983 34428
rect 57039 34372 57825 34428
rect 57881 34372 58465 34428
rect 58521 34372 59048 34428
rect 59104 34372 60326 34428
rect 60382 34372 60484 34428
rect 60540 34372 62528 34428
rect 62584 34372 62608 34428
rect 62664 34372 74216 34428
rect 74272 34372 74296 34428
rect 74352 34372 74376 34428
rect 74432 34372 74456 34428
rect 74512 34372 75028 34428
rect 964 34348 75028 34372
rect 964 34292 2044 34348
rect 2100 34292 5540 34348
rect 5596 34292 8430 34348
rect 8486 34292 11320 34348
rect 11376 34292 14210 34348
rect 14266 34292 17100 34348
rect 17156 34292 19990 34348
rect 20046 34292 22880 34348
rect 22936 34292 25770 34348
rect 25826 34292 28660 34348
rect 28716 34292 31550 34348
rect 31606 34292 34440 34348
rect 34496 34292 37330 34348
rect 37386 34292 40220 34348
rect 40276 34292 43110 34348
rect 43166 34292 46000 34348
rect 46056 34292 49008 34348
rect 49064 34292 52237 34348
rect 52293 34292 53638 34348
rect 53694 34292 53806 34348
rect 53862 34292 54550 34348
rect 54606 34292 54940 34348
rect 54996 34292 55656 34348
rect 55712 34292 56234 34348
rect 56290 34292 56679 34348
rect 56735 34292 56983 34348
rect 57039 34292 57825 34348
rect 57881 34292 58465 34348
rect 58521 34292 59048 34348
rect 59104 34292 60326 34348
rect 60382 34292 60484 34348
rect 60540 34292 62528 34348
rect 62584 34292 62608 34348
rect 62664 34292 74216 34348
rect 74272 34292 74296 34348
rect 74352 34292 74376 34348
rect 74432 34292 74456 34348
rect 74512 34292 75028 34348
rect 964 34264 75028 34292
rect 964 32236 75028 32264
rect 964 32180 2184 32236
rect 2240 32180 2264 32236
rect 2320 32180 5393 32236
rect 5449 32180 8283 32236
rect 8339 32180 11173 32236
rect 11229 32180 14063 32236
rect 14119 32180 16953 32236
rect 17009 32180 19843 32236
rect 19899 32180 22733 32236
rect 22789 32180 25623 32236
rect 25679 32180 28513 32236
rect 28569 32180 31403 32236
rect 31459 32180 34293 32236
rect 34349 32180 37183 32236
rect 37239 32180 40073 32236
rect 40129 32180 42963 32236
rect 43019 32180 45853 32236
rect 45909 32180 48800 32236
rect 48856 32180 49662 32236
rect 49718 32180 49742 32236
rect 49798 32180 52956 32236
rect 53012 32180 53114 32236
rect 53170 32180 53470 32236
rect 53526 32180 54788 32236
rect 54844 32180 55381 32236
rect 55437 32180 56527 32236
rect 56583 32180 57963 32236
rect 58019 32180 58043 32236
rect 58099 32180 59206 32236
rect 59262 32180 59364 32236
rect 59420 32180 59672 32236
rect 59728 32180 59818 32236
rect 59874 32180 59954 32236
rect 60010 32180 60034 32236
rect 60090 32180 62326 32236
rect 62382 32180 62406 32236
rect 62462 32180 71864 32236
rect 71920 32180 71944 32236
rect 72000 32180 72024 32236
rect 72080 32180 72104 32236
rect 72160 32180 75028 32236
rect 964 32156 75028 32180
rect 964 32100 2184 32156
rect 2240 32100 2264 32156
rect 2320 32100 5393 32156
rect 5449 32100 8283 32156
rect 8339 32100 11173 32156
rect 11229 32100 14063 32156
rect 14119 32100 16953 32156
rect 17009 32100 19843 32156
rect 19899 32100 22733 32156
rect 22789 32100 25623 32156
rect 25679 32100 28513 32156
rect 28569 32100 31403 32156
rect 31459 32100 34293 32156
rect 34349 32100 37183 32156
rect 37239 32100 40073 32156
rect 40129 32100 42963 32156
rect 43019 32100 45853 32156
rect 45909 32100 48800 32156
rect 48856 32100 49662 32156
rect 49718 32100 49742 32156
rect 49798 32100 52956 32156
rect 53012 32100 53114 32156
rect 53170 32100 53470 32156
rect 53526 32100 54788 32156
rect 54844 32100 55381 32156
rect 55437 32100 56527 32156
rect 56583 32100 57963 32156
rect 58019 32100 58043 32156
rect 58099 32100 59206 32156
rect 59262 32100 59364 32156
rect 59420 32100 59672 32156
rect 59728 32100 59818 32156
rect 59874 32100 59954 32156
rect 60010 32100 60034 32156
rect 60090 32100 62326 32156
rect 62382 32100 62406 32156
rect 62462 32100 71864 32156
rect 71920 32100 71944 32156
rect 72000 32100 72024 32156
rect 72080 32100 72104 32156
rect 72160 32100 75028 32156
rect 964 32076 75028 32100
rect 964 32020 2184 32076
rect 2240 32020 2264 32076
rect 2320 32020 5393 32076
rect 5449 32020 8283 32076
rect 8339 32020 11173 32076
rect 11229 32020 14063 32076
rect 14119 32020 16953 32076
rect 17009 32020 19843 32076
rect 19899 32020 22733 32076
rect 22789 32020 25623 32076
rect 25679 32020 28513 32076
rect 28569 32020 31403 32076
rect 31459 32020 34293 32076
rect 34349 32020 37183 32076
rect 37239 32020 40073 32076
rect 40129 32020 42963 32076
rect 43019 32020 45853 32076
rect 45909 32020 48800 32076
rect 48856 32020 49662 32076
rect 49718 32020 49742 32076
rect 49798 32020 52956 32076
rect 53012 32020 53114 32076
rect 53170 32020 53470 32076
rect 53526 32020 54788 32076
rect 54844 32020 55381 32076
rect 55437 32020 56527 32076
rect 56583 32020 57963 32076
rect 58019 32020 58043 32076
rect 58099 32020 59206 32076
rect 59262 32020 59364 32076
rect 59420 32020 59672 32076
rect 59728 32020 59818 32076
rect 59874 32020 59954 32076
rect 60010 32020 60034 32076
rect 60090 32020 62326 32076
rect 62382 32020 62406 32076
rect 62462 32020 71864 32076
rect 71920 32020 71944 32076
rect 72000 32020 72024 32076
rect 72080 32020 72104 32076
rect 72160 32020 75028 32076
rect 964 31996 75028 32020
rect 964 31940 2184 31996
rect 2240 31940 2264 31996
rect 2320 31940 5393 31996
rect 5449 31940 8283 31996
rect 8339 31940 11173 31996
rect 11229 31940 14063 31996
rect 14119 31940 16953 31996
rect 17009 31940 19843 31996
rect 19899 31940 22733 31996
rect 22789 31940 25623 31996
rect 25679 31940 28513 31996
rect 28569 31940 31403 31996
rect 31459 31940 34293 31996
rect 34349 31940 37183 31996
rect 37239 31940 40073 31996
rect 40129 31940 42963 31996
rect 43019 31940 45853 31996
rect 45909 31940 48800 31996
rect 48856 31940 49662 31996
rect 49718 31940 49742 31996
rect 49798 31940 52956 31996
rect 53012 31940 53114 31996
rect 53170 31940 53470 31996
rect 53526 31940 54788 31996
rect 54844 31940 55381 31996
rect 55437 31940 56527 31996
rect 56583 31940 57963 31996
rect 58019 31940 58043 31996
rect 58099 31940 59206 31996
rect 59262 31940 59364 31996
rect 59420 31940 59672 31996
rect 59728 31940 59818 31996
rect 59874 31940 59954 31996
rect 60010 31940 60034 31996
rect 60090 31940 62326 31996
rect 62382 31940 62406 31996
rect 62462 31940 71864 31996
rect 71920 31940 71944 31996
rect 72000 31940 72024 31996
rect 72080 31940 72104 31996
rect 72160 31940 75028 31996
rect 964 31912 75028 31940
rect 964 24588 75028 24616
rect 964 24532 2044 24588
rect 2100 24532 5540 24588
rect 5596 24532 8430 24588
rect 8486 24532 11320 24588
rect 11376 24532 14210 24588
rect 14266 24532 17100 24588
rect 17156 24532 19990 24588
rect 20046 24532 22880 24588
rect 22936 24532 25770 24588
rect 25826 24532 28660 24588
rect 28716 24532 31550 24588
rect 31606 24532 34440 24588
rect 34496 24532 37330 24588
rect 37386 24532 40220 24588
rect 40276 24532 43110 24588
rect 43166 24532 46000 24588
rect 46056 24532 49008 24588
rect 49064 24532 52237 24588
rect 52293 24532 53638 24588
rect 53694 24532 53806 24588
rect 53862 24532 54550 24588
rect 54606 24532 54940 24588
rect 54996 24532 55656 24588
rect 55712 24532 56234 24588
rect 56290 24532 56679 24588
rect 56735 24532 56983 24588
rect 57039 24532 57825 24588
rect 57881 24532 58465 24588
rect 58521 24532 59048 24588
rect 59104 24532 60326 24588
rect 60382 24532 60484 24588
rect 60540 24532 62528 24588
rect 62584 24532 62608 24588
rect 62664 24532 74216 24588
rect 74272 24532 74296 24588
rect 74352 24532 74376 24588
rect 74432 24532 74456 24588
rect 74512 24532 75028 24588
rect 964 24508 75028 24532
rect 964 24452 2044 24508
rect 2100 24452 5540 24508
rect 5596 24452 8430 24508
rect 8486 24452 11320 24508
rect 11376 24452 14210 24508
rect 14266 24452 17100 24508
rect 17156 24452 19990 24508
rect 20046 24452 22880 24508
rect 22936 24452 25770 24508
rect 25826 24452 28660 24508
rect 28716 24452 31550 24508
rect 31606 24452 34440 24508
rect 34496 24452 37330 24508
rect 37386 24452 40220 24508
rect 40276 24452 43110 24508
rect 43166 24452 46000 24508
rect 46056 24452 49008 24508
rect 49064 24452 52237 24508
rect 52293 24452 53638 24508
rect 53694 24452 53806 24508
rect 53862 24452 54550 24508
rect 54606 24452 54940 24508
rect 54996 24452 55656 24508
rect 55712 24452 56234 24508
rect 56290 24452 56679 24508
rect 56735 24452 56983 24508
rect 57039 24452 57825 24508
rect 57881 24452 58465 24508
rect 58521 24452 59048 24508
rect 59104 24452 60326 24508
rect 60382 24452 60484 24508
rect 60540 24452 62528 24508
rect 62584 24452 62608 24508
rect 62664 24452 74216 24508
rect 74272 24452 74296 24508
rect 74352 24452 74376 24508
rect 74432 24452 74456 24508
rect 74512 24452 75028 24508
rect 964 24428 75028 24452
rect 964 24372 2044 24428
rect 2100 24372 5540 24428
rect 5596 24372 8430 24428
rect 8486 24372 11320 24428
rect 11376 24372 14210 24428
rect 14266 24372 17100 24428
rect 17156 24372 19990 24428
rect 20046 24372 22880 24428
rect 22936 24372 25770 24428
rect 25826 24372 28660 24428
rect 28716 24372 31550 24428
rect 31606 24372 34440 24428
rect 34496 24372 37330 24428
rect 37386 24372 40220 24428
rect 40276 24372 43110 24428
rect 43166 24372 46000 24428
rect 46056 24372 49008 24428
rect 49064 24372 52237 24428
rect 52293 24372 53638 24428
rect 53694 24372 53806 24428
rect 53862 24372 54550 24428
rect 54606 24372 54940 24428
rect 54996 24372 55656 24428
rect 55712 24372 56234 24428
rect 56290 24372 56679 24428
rect 56735 24372 56983 24428
rect 57039 24372 57825 24428
rect 57881 24372 58465 24428
rect 58521 24372 59048 24428
rect 59104 24372 60326 24428
rect 60382 24372 60484 24428
rect 60540 24372 62528 24428
rect 62584 24372 62608 24428
rect 62664 24372 74216 24428
rect 74272 24372 74296 24428
rect 74352 24372 74376 24428
rect 74432 24372 74456 24428
rect 74512 24372 75028 24428
rect 964 24348 75028 24372
rect 964 24292 2044 24348
rect 2100 24292 5540 24348
rect 5596 24292 8430 24348
rect 8486 24292 11320 24348
rect 11376 24292 14210 24348
rect 14266 24292 17100 24348
rect 17156 24292 19990 24348
rect 20046 24292 22880 24348
rect 22936 24292 25770 24348
rect 25826 24292 28660 24348
rect 28716 24292 31550 24348
rect 31606 24292 34440 24348
rect 34496 24292 37330 24348
rect 37386 24292 40220 24348
rect 40276 24292 43110 24348
rect 43166 24292 46000 24348
rect 46056 24292 49008 24348
rect 49064 24292 52237 24348
rect 52293 24292 53638 24348
rect 53694 24292 53806 24348
rect 53862 24292 54550 24348
rect 54606 24292 54940 24348
rect 54996 24292 55656 24348
rect 55712 24292 56234 24348
rect 56290 24292 56679 24348
rect 56735 24292 56983 24348
rect 57039 24292 57825 24348
rect 57881 24292 58465 24348
rect 58521 24292 59048 24348
rect 59104 24292 60326 24348
rect 60382 24292 60484 24348
rect 60540 24292 62528 24348
rect 62584 24292 62608 24348
rect 62664 24292 74216 24348
rect 74272 24292 74296 24348
rect 74352 24292 74376 24348
rect 74432 24292 74456 24348
rect 74512 24292 75028 24348
rect 964 24264 75028 24292
rect 65425 23218 65491 23221
rect 65425 23216 65626 23218
rect 65425 23160 65430 23216
rect 65486 23160 65626 23216
rect 65425 23158 65626 23160
rect 65425 23155 65491 23158
rect 65566 22541 65626 23158
rect 65566 22536 65675 22541
rect 65566 22480 65614 22536
rect 65670 22480 65675 22536
rect 65566 22478 65675 22480
rect 65609 22475 65675 22478
rect 964 22236 75028 22264
rect 964 22180 2184 22236
rect 2240 22180 2264 22236
rect 2320 22180 5393 22236
rect 5449 22180 8283 22236
rect 8339 22180 11173 22236
rect 11229 22180 14063 22236
rect 14119 22180 16953 22236
rect 17009 22180 19843 22236
rect 19899 22180 22733 22236
rect 22789 22180 25623 22236
rect 25679 22180 28513 22236
rect 28569 22180 31403 22236
rect 31459 22180 34293 22236
rect 34349 22180 37183 22236
rect 37239 22180 40073 22236
rect 40129 22180 42963 22236
rect 43019 22180 45853 22236
rect 45909 22180 48800 22236
rect 48856 22180 49662 22236
rect 49718 22180 49742 22236
rect 49798 22180 52956 22236
rect 53012 22180 53114 22236
rect 53170 22180 53470 22236
rect 53526 22180 54788 22236
rect 54844 22180 55381 22236
rect 55437 22180 56527 22236
rect 56583 22180 57963 22236
rect 58019 22180 58043 22236
rect 58099 22180 59206 22236
rect 59262 22180 59364 22236
rect 59420 22180 59672 22236
rect 59728 22180 59818 22236
rect 59874 22180 59954 22236
rect 60010 22180 60034 22236
rect 60090 22180 62326 22236
rect 62382 22180 62406 22236
rect 62462 22180 71864 22236
rect 71920 22180 71944 22236
rect 72000 22180 72024 22236
rect 72080 22180 72104 22236
rect 72160 22180 75028 22236
rect 964 22156 75028 22180
rect 964 22100 2184 22156
rect 2240 22100 2264 22156
rect 2320 22100 5393 22156
rect 5449 22100 8283 22156
rect 8339 22100 11173 22156
rect 11229 22100 14063 22156
rect 14119 22100 16953 22156
rect 17009 22100 19843 22156
rect 19899 22100 22733 22156
rect 22789 22100 25623 22156
rect 25679 22100 28513 22156
rect 28569 22100 31403 22156
rect 31459 22100 34293 22156
rect 34349 22100 37183 22156
rect 37239 22100 40073 22156
rect 40129 22100 42963 22156
rect 43019 22100 45853 22156
rect 45909 22100 48800 22156
rect 48856 22100 49662 22156
rect 49718 22100 49742 22156
rect 49798 22100 52956 22156
rect 53012 22100 53114 22156
rect 53170 22100 53470 22156
rect 53526 22100 54788 22156
rect 54844 22100 55381 22156
rect 55437 22100 56527 22156
rect 56583 22100 57963 22156
rect 58019 22100 58043 22156
rect 58099 22100 59206 22156
rect 59262 22100 59364 22156
rect 59420 22100 59672 22156
rect 59728 22100 59818 22156
rect 59874 22100 59954 22156
rect 60010 22100 60034 22156
rect 60090 22100 62326 22156
rect 62382 22100 62406 22156
rect 62462 22100 71864 22156
rect 71920 22100 71944 22156
rect 72000 22100 72024 22156
rect 72080 22100 72104 22156
rect 72160 22100 75028 22156
rect 964 22076 75028 22100
rect 964 22020 2184 22076
rect 2240 22020 2264 22076
rect 2320 22020 5393 22076
rect 5449 22020 8283 22076
rect 8339 22020 11173 22076
rect 11229 22020 14063 22076
rect 14119 22020 16953 22076
rect 17009 22020 19843 22076
rect 19899 22020 22733 22076
rect 22789 22020 25623 22076
rect 25679 22020 28513 22076
rect 28569 22020 31403 22076
rect 31459 22020 34293 22076
rect 34349 22020 37183 22076
rect 37239 22020 40073 22076
rect 40129 22020 42963 22076
rect 43019 22020 45853 22076
rect 45909 22020 48800 22076
rect 48856 22020 49662 22076
rect 49718 22020 49742 22076
rect 49798 22020 52956 22076
rect 53012 22020 53114 22076
rect 53170 22020 53470 22076
rect 53526 22020 54788 22076
rect 54844 22020 55381 22076
rect 55437 22020 56527 22076
rect 56583 22020 57963 22076
rect 58019 22020 58043 22076
rect 58099 22020 59206 22076
rect 59262 22020 59364 22076
rect 59420 22020 59672 22076
rect 59728 22020 59818 22076
rect 59874 22020 59954 22076
rect 60010 22020 60034 22076
rect 60090 22020 62326 22076
rect 62382 22020 62406 22076
rect 62462 22020 71864 22076
rect 71920 22020 71944 22076
rect 72000 22020 72024 22076
rect 72080 22020 72104 22076
rect 72160 22020 75028 22076
rect 964 21996 75028 22020
rect 964 21940 2184 21996
rect 2240 21940 2264 21996
rect 2320 21940 5393 21996
rect 5449 21940 8283 21996
rect 8339 21940 11173 21996
rect 11229 21940 14063 21996
rect 14119 21940 16953 21996
rect 17009 21940 19843 21996
rect 19899 21940 22733 21996
rect 22789 21940 25623 21996
rect 25679 21940 28513 21996
rect 28569 21940 31403 21996
rect 31459 21940 34293 21996
rect 34349 21940 37183 21996
rect 37239 21940 40073 21996
rect 40129 21940 42963 21996
rect 43019 21940 45853 21996
rect 45909 21940 48800 21996
rect 48856 21940 49662 21996
rect 49718 21940 49742 21996
rect 49798 21940 52956 21996
rect 53012 21940 53114 21996
rect 53170 21940 53470 21996
rect 53526 21940 54788 21996
rect 54844 21940 55381 21996
rect 55437 21940 56527 21996
rect 56583 21940 57963 21996
rect 58019 21940 58043 21996
rect 58099 21940 59206 21996
rect 59262 21940 59364 21996
rect 59420 21940 59672 21996
rect 59728 21940 59818 21996
rect 59874 21940 59954 21996
rect 60010 21940 60034 21996
rect 60090 21940 62326 21996
rect 62382 21940 62406 21996
rect 62462 21940 71864 21996
rect 71920 21940 71944 21996
rect 72000 21940 72024 21996
rect 72080 21940 72104 21996
rect 72160 21940 75028 21996
rect 964 21912 75028 21940
rect 964 14588 75028 14616
rect 964 14532 2044 14588
rect 2100 14532 5540 14588
rect 5596 14532 8430 14588
rect 8486 14532 11320 14588
rect 11376 14532 14210 14588
rect 14266 14532 17100 14588
rect 17156 14532 19990 14588
rect 20046 14532 22880 14588
rect 22936 14532 25770 14588
rect 25826 14532 28660 14588
rect 28716 14532 31550 14588
rect 31606 14532 34440 14588
rect 34496 14532 37330 14588
rect 37386 14532 40220 14588
rect 40276 14532 43110 14588
rect 43166 14532 46000 14588
rect 46056 14532 49008 14588
rect 49064 14532 52237 14588
rect 52293 14532 53638 14588
rect 53694 14532 53806 14588
rect 53862 14532 54550 14588
rect 54606 14532 54940 14588
rect 54996 14532 55656 14588
rect 55712 14532 56234 14588
rect 56290 14532 56679 14588
rect 56735 14532 56983 14588
rect 57039 14532 57825 14588
rect 57881 14532 58465 14588
rect 58521 14532 59048 14588
rect 59104 14532 60326 14588
rect 60382 14532 60484 14588
rect 60540 14532 62528 14588
rect 62584 14532 62608 14588
rect 62664 14532 74216 14588
rect 74272 14532 74296 14588
rect 74352 14532 74376 14588
rect 74432 14532 74456 14588
rect 74512 14532 75028 14588
rect 964 14508 75028 14532
rect 964 14452 2044 14508
rect 2100 14452 5540 14508
rect 5596 14452 8430 14508
rect 8486 14452 11320 14508
rect 11376 14452 14210 14508
rect 14266 14452 17100 14508
rect 17156 14452 19990 14508
rect 20046 14452 22880 14508
rect 22936 14452 25770 14508
rect 25826 14452 28660 14508
rect 28716 14452 31550 14508
rect 31606 14452 34440 14508
rect 34496 14452 37330 14508
rect 37386 14452 40220 14508
rect 40276 14452 43110 14508
rect 43166 14452 46000 14508
rect 46056 14452 49008 14508
rect 49064 14452 52237 14508
rect 52293 14452 53638 14508
rect 53694 14452 53806 14508
rect 53862 14452 54550 14508
rect 54606 14452 54940 14508
rect 54996 14452 55656 14508
rect 55712 14452 56234 14508
rect 56290 14452 56679 14508
rect 56735 14452 56983 14508
rect 57039 14452 57825 14508
rect 57881 14452 58465 14508
rect 58521 14452 59048 14508
rect 59104 14452 60326 14508
rect 60382 14452 60484 14508
rect 60540 14452 62528 14508
rect 62584 14452 62608 14508
rect 62664 14452 74216 14508
rect 74272 14452 74296 14508
rect 74352 14452 74376 14508
rect 74432 14452 74456 14508
rect 74512 14452 75028 14508
rect 964 14428 75028 14452
rect 964 14372 2044 14428
rect 2100 14372 5540 14428
rect 5596 14372 8430 14428
rect 8486 14372 11320 14428
rect 11376 14372 14210 14428
rect 14266 14372 17100 14428
rect 17156 14372 19990 14428
rect 20046 14372 22880 14428
rect 22936 14372 25770 14428
rect 25826 14372 28660 14428
rect 28716 14372 31550 14428
rect 31606 14372 34440 14428
rect 34496 14372 37330 14428
rect 37386 14372 40220 14428
rect 40276 14372 43110 14428
rect 43166 14372 46000 14428
rect 46056 14372 49008 14428
rect 49064 14372 52237 14428
rect 52293 14372 53638 14428
rect 53694 14372 53806 14428
rect 53862 14372 54550 14428
rect 54606 14372 54940 14428
rect 54996 14372 55656 14428
rect 55712 14372 56234 14428
rect 56290 14372 56679 14428
rect 56735 14372 56983 14428
rect 57039 14372 57825 14428
rect 57881 14372 58465 14428
rect 58521 14372 59048 14428
rect 59104 14372 60326 14428
rect 60382 14372 60484 14428
rect 60540 14372 62528 14428
rect 62584 14372 62608 14428
rect 62664 14372 74216 14428
rect 74272 14372 74296 14428
rect 74352 14372 74376 14428
rect 74432 14372 74456 14428
rect 74512 14372 75028 14428
rect 964 14348 75028 14372
rect 964 14292 2044 14348
rect 2100 14292 5540 14348
rect 5596 14292 8430 14348
rect 8486 14292 11320 14348
rect 11376 14292 14210 14348
rect 14266 14292 17100 14348
rect 17156 14292 19990 14348
rect 20046 14292 22880 14348
rect 22936 14292 25770 14348
rect 25826 14292 28660 14348
rect 28716 14292 31550 14348
rect 31606 14292 34440 14348
rect 34496 14292 37330 14348
rect 37386 14292 40220 14348
rect 40276 14292 43110 14348
rect 43166 14292 46000 14348
rect 46056 14292 49008 14348
rect 49064 14292 52237 14348
rect 52293 14292 53638 14348
rect 53694 14292 53806 14348
rect 53862 14292 54550 14348
rect 54606 14292 54940 14348
rect 54996 14292 55656 14348
rect 55712 14292 56234 14348
rect 56290 14292 56679 14348
rect 56735 14292 56983 14348
rect 57039 14292 57825 14348
rect 57881 14292 58465 14348
rect 58521 14292 59048 14348
rect 59104 14292 60326 14348
rect 60382 14292 60484 14348
rect 60540 14292 62528 14348
rect 62584 14292 62608 14348
rect 62664 14292 74216 14348
rect 74272 14292 74296 14348
rect 74352 14292 74376 14348
rect 74432 14292 74456 14348
rect 74512 14292 75028 14348
rect 964 14264 75028 14292
rect 964 12236 75028 12264
rect 964 12180 2184 12236
rect 2240 12180 2264 12236
rect 2320 12180 5393 12236
rect 5449 12180 8283 12236
rect 8339 12180 11173 12236
rect 11229 12180 14063 12236
rect 14119 12180 16953 12236
rect 17009 12180 19843 12236
rect 19899 12180 22733 12236
rect 22789 12180 25623 12236
rect 25679 12180 28513 12236
rect 28569 12180 31403 12236
rect 31459 12180 34293 12236
rect 34349 12180 37183 12236
rect 37239 12180 40073 12236
rect 40129 12180 42963 12236
rect 43019 12180 45853 12236
rect 45909 12180 48800 12236
rect 48856 12180 49662 12236
rect 49718 12180 49742 12236
rect 49798 12180 52956 12236
rect 53012 12180 53114 12236
rect 53170 12180 53470 12236
rect 53526 12180 54788 12236
rect 54844 12180 55381 12236
rect 55437 12180 56527 12236
rect 56583 12180 57963 12236
rect 58019 12180 58043 12236
rect 58099 12180 59206 12236
rect 59262 12180 59364 12236
rect 59420 12180 59672 12236
rect 59728 12180 59818 12236
rect 59874 12180 59954 12236
rect 60010 12180 60034 12236
rect 60090 12180 62326 12236
rect 62382 12180 62406 12236
rect 62462 12180 71864 12236
rect 71920 12180 71944 12236
rect 72000 12180 72024 12236
rect 72080 12180 72104 12236
rect 72160 12180 75028 12236
rect 964 12156 75028 12180
rect 964 12100 2184 12156
rect 2240 12100 2264 12156
rect 2320 12100 5393 12156
rect 5449 12100 8283 12156
rect 8339 12100 11173 12156
rect 11229 12100 14063 12156
rect 14119 12100 16953 12156
rect 17009 12100 19843 12156
rect 19899 12100 22733 12156
rect 22789 12100 25623 12156
rect 25679 12100 28513 12156
rect 28569 12100 31403 12156
rect 31459 12100 34293 12156
rect 34349 12100 37183 12156
rect 37239 12100 40073 12156
rect 40129 12100 42963 12156
rect 43019 12100 45853 12156
rect 45909 12100 48800 12156
rect 48856 12100 49662 12156
rect 49718 12100 49742 12156
rect 49798 12100 52956 12156
rect 53012 12100 53114 12156
rect 53170 12100 53470 12156
rect 53526 12100 54788 12156
rect 54844 12100 55381 12156
rect 55437 12100 56527 12156
rect 56583 12100 57963 12156
rect 58019 12100 58043 12156
rect 58099 12100 59206 12156
rect 59262 12100 59364 12156
rect 59420 12100 59672 12156
rect 59728 12100 59818 12156
rect 59874 12100 59954 12156
rect 60010 12100 60034 12156
rect 60090 12100 62326 12156
rect 62382 12100 62406 12156
rect 62462 12100 71864 12156
rect 71920 12100 71944 12156
rect 72000 12100 72024 12156
rect 72080 12100 72104 12156
rect 72160 12100 75028 12156
rect 964 12076 75028 12100
rect 964 12020 2184 12076
rect 2240 12020 2264 12076
rect 2320 12020 5393 12076
rect 5449 12020 8283 12076
rect 8339 12020 11173 12076
rect 11229 12020 14063 12076
rect 14119 12020 16953 12076
rect 17009 12020 19843 12076
rect 19899 12020 22733 12076
rect 22789 12020 25623 12076
rect 25679 12020 28513 12076
rect 28569 12020 31403 12076
rect 31459 12020 34293 12076
rect 34349 12020 37183 12076
rect 37239 12020 40073 12076
rect 40129 12020 42963 12076
rect 43019 12020 45853 12076
rect 45909 12020 48800 12076
rect 48856 12020 49662 12076
rect 49718 12020 49742 12076
rect 49798 12020 52956 12076
rect 53012 12020 53114 12076
rect 53170 12020 53470 12076
rect 53526 12020 54788 12076
rect 54844 12020 55381 12076
rect 55437 12020 56527 12076
rect 56583 12020 57963 12076
rect 58019 12020 58043 12076
rect 58099 12020 59206 12076
rect 59262 12020 59364 12076
rect 59420 12020 59672 12076
rect 59728 12020 59818 12076
rect 59874 12020 59954 12076
rect 60010 12020 60034 12076
rect 60090 12020 62326 12076
rect 62382 12020 62406 12076
rect 62462 12020 71864 12076
rect 71920 12020 71944 12076
rect 72000 12020 72024 12076
rect 72080 12020 72104 12076
rect 72160 12020 75028 12076
rect 964 11996 75028 12020
rect 964 11940 2184 11996
rect 2240 11940 2264 11996
rect 2320 11940 5393 11996
rect 5449 11940 8283 11996
rect 8339 11940 11173 11996
rect 11229 11940 14063 11996
rect 14119 11940 16953 11996
rect 17009 11940 19843 11996
rect 19899 11940 22733 11996
rect 22789 11940 25623 11996
rect 25679 11940 28513 11996
rect 28569 11940 31403 11996
rect 31459 11940 34293 11996
rect 34349 11940 37183 11996
rect 37239 11940 40073 11996
rect 40129 11940 42963 11996
rect 43019 11940 45853 11996
rect 45909 11940 48800 11996
rect 48856 11940 49662 11996
rect 49718 11940 49742 11996
rect 49798 11940 52956 11996
rect 53012 11940 53114 11996
rect 53170 11940 53470 11996
rect 53526 11940 54788 11996
rect 54844 11940 55381 11996
rect 55437 11940 56527 11996
rect 56583 11940 57963 11996
rect 58019 11940 58043 11996
rect 58099 11940 59206 11996
rect 59262 11940 59364 11996
rect 59420 11940 59672 11996
rect 59728 11940 59818 11996
rect 59874 11940 59954 11996
rect 60010 11940 60034 11996
rect 60090 11940 62326 11996
rect 62382 11940 62406 11996
rect 62462 11940 71864 11996
rect 71920 11940 71944 11996
rect 72000 11940 72024 11996
rect 72080 11940 72104 11996
rect 72160 11940 75028 11996
rect 964 11912 75028 11940
rect 64873 7986 64939 7989
rect 64873 7984 65258 7986
rect 64873 7928 64878 7984
rect 64934 7928 65258 7984
rect 64873 7926 65258 7928
rect 64873 7923 64939 7926
rect 65198 7445 65258 7926
rect 65198 7440 65307 7445
rect 65198 7384 65246 7440
rect 65302 7384 65307 7440
rect 65198 7382 65307 7384
rect 65241 7379 65307 7382
rect 60917 6626 60983 6629
rect 61377 6626 61443 6629
rect 60917 6624 61443 6626
rect 60917 6568 60922 6624
rect 60978 6568 61382 6624
rect 61438 6568 61443 6624
rect 60917 6566 61443 6568
rect 60917 6563 60983 6566
rect 61377 6563 61443 6566
rect 58525 6354 58591 6357
rect 65793 6354 65859 6357
rect 58525 6352 65859 6354
rect 58525 6296 58530 6352
rect 58586 6296 65798 6352
rect 65854 6296 65859 6352
rect 58525 6294 65859 6296
rect 58525 6291 58591 6294
rect 65793 6291 65859 6294
rect 57605 6218 57671 6221
rect 71313 6218 71379 6221
rect 57605 6216 71379 6218
rect 57605 6160 57610 6216
rect 57666 6160 71318 6216
rect 71374 6160 71379 6216
rect 57605 6158 71379 6160
rect 57605 6155 57671 6158
rect 71313 6155 71379 6158
rect 41689 6082 41755 6085
rect 64137 6082 64203 6085
rect 64413 6082 64479 6085
rect 41689 6080 64203 6082
rect 41689 6024 41694 6080
rect 41750 6024 64142 6080
rect 64198 6024 64203 6080
rect 41689 6022 64203 6024
rect 41689 6019 41755 6022
rect 64137 6019 64203 6022
rect 64278 6080 64479 6082
rect 64278 6024 64418 6080
rect 64474 6024 64479 6080
rect 64278 6022 64479 6024
rect 39481 5946 39547 5949
rect 62665 5946 62731 5949
rect 39481 5944 62731 5946
rect 39481 5888 39486 5944
rect 39542 5888 62670 5944
rect 62726 5888 62731 5944
rect 39481 5886 62731 5888
rect 39481 5883 39547 5886
rect 62665 5883 62731 5886
rect 40401 5810 40467 5813
rect 64278 5810 64338 6022
rect 64413 6019 64479 6022
rect 40401 5808 64338 5810
rect 40401 5752 40406 5808
rect 40462 5752 64338 5808
rect 40401 5750 64338 5752
rect 40401 5747 40467 5750
rect 38745 5674 38811 5677
rect 66621 5674 66687 5677
rect 38745 5672 66687 5674
rect 38745 5616 38750 5672
rect 38806 5616 66626 5672
rect 66682 5616 66687 5672
rect 38745 5614 66687 5616
rect 38745 5611 38811 5614
rect 66621 5611 66687 5614
rect 44081 5266 44147 5269
rect 46197 5266 46263 5269
rect 44081 5264 46263 5266
rect 44081 5208 44086 5264
rect 44142 5208 46202 5264
rect 46258 5208 46263 5264
rect 44081 5206 46263 5208
rect 44081 5203 44147 5206
rect 46197 5203 46263 5206
rect 52821 5266 52887 5269
rect 56593 5266 56659 5269
rect 52821 5264 56659 5266
rect 52821 5208 52826 5264
rect 52882 5208 56598 5264
rect 56654 5208 56659 5264
rect 52821 5206 56659 5208
rect 52821 5203 52887 5206
rect 56593 5203 56659 5206
rect 39205 5130 39271 5133
rect 46657 5130 46723 5133
rect 39205 5128 46723 5130
rect 39205 5072 39210 5128
rect 39266 5072 46662 5128
rect 46718 5072 46723 5128
rect 39205 5070 46723 5072
rect 39205 5067 39271 5070
rect 46657 5067 46723 5070
rect 51257 5130 51323 5133
rect 54845 5130 54911 5133
rect 51257 5128 54911 5130
rect 51257 5072 51262 5128
rect 51318 5072 54850 5128
rect 54906 5072 54911 5128
rect 51257 5070 54911 5072
rect 51257 5067 51323 5070
rect 54845 5067 54911 5070
rect 40585 4858 40651 4861
rect 47577 4858 47643 4861
rect 40585 4856 47643 4858
rect 40585 4800 40590 4856
rect 40646 4800 47582 4856
rect 47638 4800 47643 4856
rect 40585 4798 47643 4800
rect 40585 4795 40651 4798
rect 47577 4795 47643 4798
rect 964 4588 75028 4616
rect 964 4532 4216 4588
rect 4272 4532 4296 4588
rect 4352 4532 4376 4588
rect 4432 4532 4456 4588
rect 4512 4532 14216 4588
rect 14272 4532 14296 4588
rect 14352 4532 14376 4588
rect 14432 4532 14456 4588
rect 14512 4532 24216 4588
rect 24272 4532 24296 4588
rect 24352 4532 24376 4588
rect 24432 4532 24456 4588
rect 24512 4532 34216 4588
rect 34272 4532 34296 4588
rect 34352 4532 34376 4588
rect 34432 4532 34456 4588
rect 34512 4532 44216 4588
rect 44272 4532 44296 4588
rect 44352 4532 44376 4588
rect 44432 4532 44456 4588
rect 44512 4532 54216 4588
rect 54272 4532 54296 4588
rect 54352 4532 54376 4588
rect 54432 4532 54456 4588
rect 54512 4532 64216 4588
rect 64272 4532 64296 4588
rect 64352 4532 64376 4588
rect 64432 4532 64456 4588
rect 64512 4532 74216 4588
rect 74272 4532 74296 4588
rect 74352 4532 74376 4588
rect 74432 4532 74456 4588
rect 74512 4532 75028 4588
rect 964 4508 75028 4532
rect 964 4452 4216 4508
rect 4272 4452 4296 4508
rect 4352 4452 4376 4508
rect 4432 4452 4456 4508
rect 4512 4452 14216 4508
rect 14272 4452 14296 4508
rect 14352 4452 14376 4508
rect 14432 4452 14456 4508
rect 14512 4452 24216 4508
rect 24272 4452 24296 4508
rect 24352 4452 24376 4508
rect 24432 4452 24456 4508
rect 24512 4452 34216 4508
rect 34272 4452 34296 4508
rect 34352 4452 34376 4508
rect 34432 4452 34456 4508
rect 34512 4452 44216 4508
rect 44272 4452 44296 4508
rect 44352 4452 44376 4508
rect 44432 4452 44456 4508
rect 44512 4452 54216 4508
rect 54272 4452 54296 4508
rect 54352 4452 54376 4508
rect 54432 4452 54456 4508
rect 54512 4452 64216 4508
rect 64272 4452 64296 4508
rect 64352 4452 64376 4508
rect 64432 4452 64456 4508
rect 64512 4452 74216 4508
rect 74272 4452 74296 4508
rect 74352 4452 74376 4508
rect 74432 4452 74456 4508
rect 74512 4452 75028 4508
rect 964 4428 75028 4452
rect 964 4372 4216 4428
rect 4272 4372 4296 4428
rect 4352 4372 4376 4428
rect 4432 4372 4456 4428
rect 4512 4372 14216 4428
rect 14272 4372 14296 4428
rect 14352 4372 14376 4428
rect 14432 4372 14456 4428
rect 14512 4372 24216 4428
rect 24272 4372 24296 4428
rect 24352 4372 24376 4428
rect 24432 4372 24456 4428
rect 24512 4372 34216 4428
rect 34272 4372 34296 4428
rect 34352 4372 34376 4428
rect 34432 4372 34456 4428
rect 34512 4372 44216 4428
rect 44272 4372 44296 4428
rect 44352 4372 44376 4428
rect 44432 4372 44456 4428
rect 44512 4372 54216 4428
rect 54272 4372 54296 4428
rect 54352 4372 54376 4428
rect 54432 4372 54456 4428
rect 54512 4372 64216 4428
rect 64272 4372 64296 4428
rect 64352 4372 64376 4428
rect 64432 4372 64456 4428
rect 64512 4372 74216 4428
rect 74272 4372 74296 4428
rect 74352 4372 74376 4428
rect 74432 4372 74456 4428
rect 74512 4372 75028 4428
rect 964 4348 75028 4372
rect 964 4292 4216 4348
rect 4272 4292 4296 4348
rect 4352 4292 4376 4348
rect 4432 4292 4456 4348
rect 4512 4292 14216 4348
rect 14272 4292 14296 4348
rect 14352 4292 14376 4348
rect 14432 4292 14456 4348
rect 14512 4292 24216 4348
rect 24272 4292 24296 4348
rect 24352 4292 24376 4348
rect 24432 4292 24456 4348
rect 24512 4292 34216 4348
rect 34272 4292 34296 4348
rect 34352 4292 34376 4348
rect 34432 4292 34456 4348
rect 34512 4292 44216 4348
rect 44272 4292 44296 4348
rect 44352 4292 44376 4348
rect 44432 4292 44456 4348
rect 44512 4292 54216 4348
rect 54272 4292 54296 4348
rect 54352 4292 54376 4348
rect 54432 4292 54456 4348
rect 54512 4292 64216 4348
rect 64272 4292 64296 4348
rect 64352 4292 64376 4348
rect 64432 4292 64456 4348
rect 64512 4292 74216 4348
rect 74272 4292 74296 4348
rect 74352 4292 74376 4348
rect 74432 4292 74456 4348
rect 74512 4292 75028 4348
rect 964 4264 75028 4292
rect 41321 4042 41387 4045
rect 44081 4042 44147 4045
rect 41321 4040 44147 4042
rect 41321 3984 41326 4040
rect 41382 3984 44086 4040
rect 44142 3984 44147 4040
rect 41321 3982 44147 3984
rect 41321 3979 41387 3982
rect 44081 3979 44147 3982
rect 40861 3770 40927 3773
rect 47853 3770 47919 3773
rect 40861 3768 47919 3770
rect 40861 3712 40866 3768
rect 40922 3712 47858 3768
rect 47914 3712 47919 3768
rect 40861 3710 47919 3712
rect 40861 3707 40927 3710
rect 47853 3707 47919 3710
rect 40309 3634 40375 3637
rect 45093 3634 45159 3637
rect 40309 3632 45159 3634
rect 40309 3576 40314 3632
rect 40370 3576 45098 3632
rect 45154 3576 45159 3632
rect 40309 3574 45159 3576
rect 40309 3571 40375 3574
rect 45093 3571 45159 3574
rect 23013 3362 23079 3365
rect 69013 3362 69079 3365
rect 23013 3360 69079 3362
rect 23013 3304 23018 3360
rect 23074 3304 69018 3360
rect 69074 3304 69079 3360
rect 23013 3302 69079 3304
rect 23013 3299 23079 3302
rect 69013 3299 69079 3302
rect 42333 3090 42399 3093
rect 47945 3090 48011 3093
rect 42333 3088 48011 3090
rect 42333 3032 42338 3088
rect 42394 3032 47950 3088
rect 48006 3032 48011 3088
rect 42333 3030 48011 3032
rect 42333 3027 42399 3030
rect 47945 3027 48011 3030
rect 41689 2954 41755 2957
rect 42701 2954 42767 2957
rect 41689 2952 42767 2954
rect 41689 2896 41694 2952
rect 41750 2896 42706 2952
rect 42762 2896 42767 2952
rect 41689 2894 42767 2896
rect 41689 2891 41755 2894
rect 42701 2891 42767 2894
rect 964 2236 75028 2264
rect 964 2180 1864 2236
rect 1920 2180 1944 2236
rect 2000 2180 2024 2236
rect 2080 2180 2104 2236
rect 2160 2180 11864 2236
rect 11920 2180 11944 2236
rect 12000 2180 12024 2236
rect 12080 2180 12104 2236
rect 12160 2180 21864 2236
rect 21920 2180 21944 2236
rect 22000 2180 22024 2236
rect 22080 2180 22104 2236
rect 22160 2180 31864 2236
rect 31920 2180 31944 2236
rect 32000 2180 32024 2236
rect 32080 2180 32104 2236
rect 32160 2180 41864 2236
rect 41920 2180 41944 2236
rect 42000 2180 42024 2236
rect 42080 2180 42104 2236
rect 42160 2180 51864 2236
rect 51920 2180 51944 2236
rect 52000 2180 52024 2236
rect 52080 2180 52104 2236
rect 52160 2180 61864 2236
rect 61920 2180 61944 2236
rect 62000 2180 62024 2236
rect 62080 2180 62104 2236
rect 62160 2180 71864 2236
rect 71920 2180 71944 2236
rect 72000 2180 72024 2236
rect 72080 2180 72104 2236
rect 72160 2180 75028 2236
rect 964 2156 75028 2180
rect 964 2100 1864 2156
rect 1920 2100 1944 2156
rect 2000 2100 2024 2156
rect 2080 2100 2104 2156
rect 2160 2100 11864 2156
rect 11920 2100 11944 2156
rect 12000 2100 12024 2156
rect 12080 2100 12104 2156
rect 12160 2100 21864 2156
rect 21920 2100 21944 2156
rect 22000 2100 22024 2156
rect 22080 2100 22104 2156
rect 22160 2100 31864 2156
rect 31920 2100 31944 2156
rect 32000 2100 32024 2156
rect 32080 2100 32104 2156
rect 32160 2100 41864 2156
rect 41920 2100 41944 2156
rect 42000 2100 42024 2156
rect 42080 2100 42104 2156
rect 42160 2100 51864 2156
rect 51920 2100 51944 2156
rect 52000 2100 52024 2156
rect 52080 2100 52104 2156
rect 52160 2100 61864 2156
rect 61920 2100 61944 2156
rect 62000 2100 62024 2156
rect 62080 2100 62104 2156
rect 62160 2100 71864 2156
rect 71920 2100 71944 2156
rect 72000 2100 72024 2156
rect 72080 2100 72104 2156
rect 72160 2100 75028 2156
rect 964 2076 75028 2100
rect 964 2020 1864 2076
rect 1920 2020 1944 2076
rect 2000 2020 2024 2076
rect 2080 2020 2104 2076
rect 2160 2020 11864 2076
rect 11920 2020 11944 2076
rect 12000 2020 12024 2076
rect 12080 2020 12104 2076
rect 12160 2020 21864 2076
rect 21920 2020 21944 2076
rect 22000 2020 22024 2076
rect 22080 2020 22104 2076
rect 22160 2020 31864 2076
rect 31920 2020 31944 2076
rect 32000 2020 32024 2076
rect 32080 2020 32104 2076
rect 32160 2020 41864 2076
rect 41920 2020 41944 2076
rect 42000 2020 42024 2076
rect 42080 2020 42104 2076
rect 42160 2020 51864 2076
rect 51920 2020 51944 2076
rect 52000 2020 52024 2076
rect 52080 2020 52104 2076
rect 52160 2020 61864 2076
rect 61920 2020 61944 2076
rect 62000 2020 62024 2076
rect 62080 2020 62104 2076
rect 62160 2020 71864 2076
rect 71920 2020 71944 2076
rect 72000 2020 72024 2076
rect 72080 2020 72104 2076
rect 72160 2020 75028 2076
rect 964 1996 75028 2020
rect 964 1940 1864 1996
rect 1920 1940 1944 1996
rect 2000 1940 2024 1996
rect 2080 1940 2104 1996
rect 2160 1940 11864 1996
rect 11920 1940 11944 1996
rect 12000 1940 12024 1996
rect 12080 1940 12104 1996
rect 12160 1940 21864 1996
rect 21920 1940 21944 1996
rect 22000 1940 22024 1996
rect 22080 1940 22104 1996
rect 22160 1940 31864 1996
rect 31920 1940 31944 1996
rect 32000 1940 32024 1996
rect 32080 1940 32104 1996
rect 32160 1940 41864 1996
rect 41920 1940 41944 1996
rect 42000 1940 42024 1996
rect 42080 1940 42104 1996
rect 42160 1940 51864 1996
rect 51920 1940 51944 1996
rect 52000 1940 52024 1996
rect 52080 1940 52104 1996
rect 52160 1940 61864 1996
rect 61920 1940 61944 1996
rect 62000 1940 62024 1996
rect 62080 1940 62104 1996
rect 62160 1940 71864 1996
rect 71920 1940 71944 1996
rect 72000 1940 72024 1996
rect 72080 1940 72104 1996
rect 72160 1940 75028 1996
rect 964 1912 75028 1940
use sky130_fd_sc_hd__clkinv_4  _13_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 33856 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _14_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 28888 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _15_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 36432 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _16_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 30084 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _17_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 28244 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _18_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 26864 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _19_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 29624 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 65964 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1704896540
transform -1 0 66700 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 65596 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_wb_clk_i
timestamp 1704896540
transform -1 0 44160 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_wb_clk_i
timestamp 1704896540
transform 1 0 65596 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__clkinv_16  clkload0 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 44528 0 1 5440
box -38 -48 2246 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1288 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1704896540
transform 1 0 2392 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3496 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1704896540
transform 1 0 3680 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1704896540
transform 1 0 4784 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5888 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1704896540
transform 1 0 6256 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1704896540
transform 1 0 7360 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1704896540
transform 1 0 8464 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1704896540
transform 1 0 8832 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1704896540
transform 1 0 9936 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1704896540
transform 1 0 11040 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1704896540
transform 1 0 11408 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1704896540
transform 1 0 12512 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1704896540
transform 1 0 13616 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1704896540
transform 1 0 13984 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1704896540
transform 1 0 15088 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 1704896540
transform 1 0 16192 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1704896540
transform 1 0 16560 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 1704896540
transform 1 0 17664 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 1704896540
transform 1 0 18768 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_197 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 19136 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_205
timestamp 1704896540
transform 1 0 19872 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_253
timestamp 1704896540
transform 1 0 24288 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_281
timestamp 1704896540
transform 1 0 26864 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_309
timestamp 1704896540
transform 1 0 29440 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_361
timestamp 1704896540
transform 1 0 34224 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_365 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 34592 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_391
timestamp 1704896540
transform 1 0 36984 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_393
timestamp 1704896540
transform 1 0 37168 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_445
timestamp 1704896540
transform 1 0 41952 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_473
timestamp 1704896540
transform 1 0 44528 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_477
timestamp 1704896540
transform 1 0 44896 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_529
timestamp 1704896540
transform 1 0 49680 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_557
timestamp 1704896540
transform 1 0 52256 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_585
timestamp 1704896540
transform 1 0 54832 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_613
timestamp 1704896540
transform 1 0 57408 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_641
timestamp 1704896540
transform 1 0 59984 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_669
timestamp 1704896540
transform 1 0 62560 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_697
timestamp 1704896540
transform 1 0 65136 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_701 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 65504 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_727
timestamp 1704896540
transform 1 0 67896 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_753
timestamp 1704896540
transform 1 0 70288 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_781
timestamp 1704896540
transform 1 0 72864 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1704896540
transform 1 0 1288 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1704896540
transform 1 0 2392 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1704896540
transform 1 0 3496 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1704896540
transform 1 0 4600 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1704896540
transform 1 0 5704 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1704896540
transform 1 0 6072 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1704896540
transform 1 0 6256 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1704896540
transform 1 0 7360 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1704896540
transform 1 0 8464 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1704896540
transform 1 0 9568 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10672 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1704896540
transform 1 0 11224 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1704896540
transform 1 0 11408 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1704896540
transform 1 0 12512 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1704896540
transform 1 0 13616 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1704896540
transform 1 0 14720 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1704896540
transform 1 0 15824 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1704896540
transform 1 0 16376 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1704896540
transform 1 0 16560 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1704896540
transform 1 0 17664 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1704896540
transform 1 0 18768 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_205
timestamp 1704896540
transform 1 0 19872 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_213
timestamp 1704896540
transform 1 0 20608 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_225
timestamp 1704896540
transform 1 0 21712 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_284
timestamp 1704896540
transform 1 0 27140 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_301
timestamp 1704896540
transform 1 0 28704 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_337
timestamp 1704896540
transform 1 0 32016 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_356
timestamp 1704896540
transform 1 0 33764 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_409
timestamp 1704896540
transform 1 0 38640 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_445
timestamp 1704896540
transform 1 0 41952 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_449
timestamp 1704896540
transform 1 0 42320 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_502
timestamp 1704896540
transform 1 0 47196 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_509
timestamp 1704896540
transform 1 0 47840 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_556
timestamp 1704896540
transform 1 0 52164 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_569
timestamp 1704896540
transform 1 0 53360 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_625
timestamp 1704896540
transform 1 0 58512 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_629
timestamp 1704896540
transform 1 0 58880 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_670
timestamp 1704896540
transform 1 0 62652 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_673
timestamp 1704896540
transform 1 0 62928 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_723
timestamp 1704896540
transform 1 0 67528 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_727
timestamp 1704896540
transform 1 0 67896 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_781
timestamp 1704896540
transform 1 0 72864 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_791
timestamp 1704896540
transform 1 0 73784 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_799
timestamp 1704896540
transform 1 0 74520 0 -1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1704896540
transform 1 0 1288 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1704896540
transform 1 0 2392 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1704896540
transform 1 0 3496 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1704896540
transform 1 0 3680 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1704896540
transform 1 0 4784 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1704896540
transform 1 0 5888 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1704896540
transform 1 0 6992 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1704896540
transform 1 0 8096 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1704896540
transform 1 0 8648 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1704896540
transform 1 0 8832 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1704896540
transform 1 0 9936 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1704896540
transform 1 0 11040 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1704896540
transform 1 0 12144 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1704896540
transform 1 0 13248 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1704896540
transform 1 0 13800 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1704896540
transform 1 0 13984 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1704896540
transform 1 0 15088 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1704896540
transform 1 0 16192 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1704896540
transform 1 0 17296 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1704896540
transform 1 0 18400 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1704896540
transform 1 0 18952 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1704896540
transform 1 0 19136 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1704896540
transform 1 0 20240 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_221
timestamp 1704896540
transform 1 0 21344 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_227
timestamp 1704896540
transform 1 0 21896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_299
timestamp 1704896540
transform 1 0 28520 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_365
timestamp 1704896540
transform 1 0 34592 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_407
timestamp 1704896540
transform 1 0 38456 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_418
timestamp 1704896540
transform 1 0 39468 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_475
timestamp 1704896540
transform 1 0 44712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_529
timestamp 1704896540
transform 1 0 49680 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_587
timestamp 1704896540
transform 1 0 55016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_643
timestamp 1704896540
transform 1 0 60168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_685
timestamp 1704896540
transform 1 0 64032 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_697
timestamp 1704896540
transform 1 0 65136 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_755
timestamp 1704896540
transform 1 0 70472 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_781
timestamp 1704896540
transform 1 0 72864 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_793
timestamp 1704896540
transform 1 0 73968 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1704896540
transform 1 0 1288 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1704896540
transform 1 0 2392 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1704896540
transform 1 0 3496 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1704896540
transform 1 0 4600 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1704896540
transform 1 0 5704 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1704896540
transform 1 0 6072 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1704896540
transform 1 0 6256 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1704896540
transform 1 0 7360 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1704896540
transform 1 0 8464 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1704896540
transform 1 0 9568 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1704896540
transform 1 0 10672 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1704896540
transform 1 0 11224 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1704896540
transform 1 0 11408 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1704896540
transform 1 0 12512 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1704896540
transform 1 0 13616 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1704896540
transform 1 0 14720 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1704896540
transform 1 0 15824 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1704896540
transform 1 0 16376 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1704896540
transform 1 0 16560 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1704896540
transform 1 0 17664 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1704896540
transform 1 0 18768 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1704896540
transform 1 0 19872 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1704896540
transform 1 0 20976 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1704896540
transform 1 0 21528 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_225
timestamp 1704896540
transform 1 0 21712 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_231
timestamp 1704896540
transform 1 0 22264 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_281
timestamp 1704896540
transform 1 0 26864 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_311
timestamp 1704896540
transform 1 0 29624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_391
timestamp 1704896540
transform 1 0 36984 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_393
timestamp 1704896540
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_424
timestamp 1704896540
transform 1 0 40020 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_441
timestamp 1704896540
transform 1 0 41584 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_501
timestamp 1704896540
transform 1 0 47104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_559
timestamp 1704896540
transform 1 0 52440 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_615
timestamp 1704896540
transform 1 0 57592 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_671
timestamp 1704896540
transform 1 0 62744 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_673
timestamp 1704896540
transform 1 0 62928 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_699
timestamp 1704896540
transform 1 0 65320 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_726
timestamp 1704896540
transform 1 0 67804 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_735
timestamp 1704896540
transform 1 0 68632 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_762
timestamp 1704896540
transform 1 0 71116 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_771
timestamp 1704896540
transform 1 0 71944 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_783
timestamp 1704896540
transform 1 0 73048 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_785
timestamp 1704896540
transform 1 0 73232 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_797
timestamp 1704896540
transform 1 0 74336 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1704896540
transform 1 0 1288 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1704896540
transform 1 0 2392 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1704896540
transform 1 0 3496 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1704896540
transform 1 0 3680 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1704896540
transform 1 0 4784 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1704896540
transform 1 0 5888 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1704896540
transform 1 0 6992 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1704896540
transform 1 0 8096 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1704896540
transform 1 0 8648 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1704896540
transform 1 0 8832 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1704896540
transform 1 0 9936 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1704896540
transform 1 0 11040 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1704896540
transform 1 0 12144 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1704896540
transform 1 0 13248 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1704896540
transform 1 0 13800 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1704896540
transform 1 0 13984 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1704896540
transform 1 0 15088 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1704896540
transform 1 0 16192 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1704896540
transform 1 0 17296 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1704896540
transform 1 0 18400 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1704896540
transform 1 0 18952 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1704896540
transform 1 0 19136 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1704896540
transform 1 0 20240 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1704896540
transform 1 0 21344 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_233
timestamp 1704896540
transform 1 0 22448 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_241
timestamp 1704896540
transform 1 0 23184 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_253
timestamp 1704896540
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_309
timestamp 1704896540
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_365
timestamp 1704896540
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_398
timestamp 1704896540
transform 1 0 37628 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_408
timestamp 1704896540
transform 1 0 38548 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_415
timestamp 1704896540
transform 1 0 39192 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_419
timestamp 1704896540
transform 1 0 39560 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_421
timestamp 1704896540
transform 1 0 39744 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_475
timestamp 1704896540
transform 1 0 44712 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_529
timestamp 1704896540
transform 1 0 49680 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_549
timestamp 1704896540
transform 1 0 51520 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_566
timestamp 1704896540
transform 1 0 53084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_578
timestamp 1704896540
transform 1 0 54188 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_586
timestamp 1704896540
transform 1 0 54924 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_597
timestamp 1704896540
transform 1 0 55936 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_609
timestamp 1704896540
transform 1 0 57040 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_613
timestamp 1704896540
transform 1 0 57408 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_628
timestamp 1704896540
transform 1 0 58788 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_640
timestamp 1704896540
transform 1 0 59892 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_645
timestamp 1704896540
transform 1 0 60352 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_652
timestamp 1704896540
transform 1 0 60996 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_664
timestamp 1704896540
transform 1 0 62100 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_676
timestamp 1704896540
transform 1 0 63204 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_684
timestamp 1704896540
transform 1 0 63940 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_691
timestamp 1704896540
transform 1 0 64584 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_699
timestamp 1704896540
transform 1 0 65320 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_701
timestamp 1704896540
transform 1 0 65504 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_713
timestamp 1704896540
transform 1 0 66608 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_725
timestamp 1704896540
transform 1 0 67712 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_737
timestamp 1704896540
transform 1 0 68816 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_749
timestamp 1704896540
transform 1 0 69920 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_755
timestamp 1704896540
transform 1 0 70472 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_757
timestamp 1704896540
transform 1 0 70656 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_769
timestamp 1704896540
transform 1 0 71760 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_781
timestamp 1704896540
transform 1 0 72864 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_793
timestamp 1704896540
transform 1 0 73968 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1704896540
transform 1 0 1288 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1704896540
transform 1 0 2392 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1704896540
transform 1 0 3496 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1704896540
transform 1 0 4600 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1704896540
transform 1 0 5704 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1704896540
transform 1 0 6072 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1704896540
transform 1 0 6256 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1704896540
transform 1 0 7360 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1704896540
transform 1 0 8464 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1704896540
transform 1 0 9568 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1704896540
transform 1 0 10672 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1704896540
transform 1 0 11224 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1704896540
transform 1 0 11408 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1704896540
transform 1 0 12512 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1704896540
transform 1 0 13616 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1704896540
transform 1 0 14720 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1704896540
transform 1 0 15824 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1704896540
transform 1 0 16376 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1704896540
transform 1 0 16560 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1704896540
transform 1 0 17664 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1704896540
transform 1 0 18768 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1704896540
transform 1 0 19872 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1704896540
transform 1 0 20976 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1704896540
transform 1 0 21528 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1704896540
transform 1 0 21712 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1704896540
transform 1 0 22816 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_249
timestamp 1704896540
transform 1 0 23920 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_255
timestamp 1704896540
transform 1 0 24472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_327
timestamp 1704896540
transform 1 0 31096 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_345
timestamp 1704896540
transform 1 0 32752 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_378
timestamp 1704896540
transform 1 0 35788 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_388
timestamp 1704896540
transform 1 0 36708 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_393
timestamp 1704896540
transform 1 0 37168 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_401
timestamp 1704896540
transform 1 0 37904 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_413
timestamp 1704896540
transform 1 0 39008 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_425
timestamp 1704896540
transform 1 0 40112 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_437
timestamp 1704896540
transform 1 0 41216 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_457
timestamp 1704896540
transform 1 0 43056 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_469
timestamp 1704896540
transform 1 0 44160 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_478
timestamp 1704896540
transform 1 0 44988 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_482
timestamp 1704896540
transform 1 0 45356 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_491
timestamp 1704896540
transform 1 0 46184 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_503
timestamp 1704896540
transform 1 0 47288 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_505
timestamp 1704896540
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_514
timestamp 1704896540
transform 1 0 48300 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_526
timestamp 1704896540
transform 1 0 49404 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_538
timestamp 1704896540
transform 1 0 50508 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_550
timestamp 1704896540
transform 1 0 51612 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_558
timestamp 1704896540
transform 1 0 52348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_561
timestamp 1704896540
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_570
timestamp 1704896540
transform 1 0 53452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_582
timestamp 1704896540
transform 1 0 54556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_594
timestamp 1704896540
transform 1 0 55660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_606
timestamp 1704896540
transform 1 0 56764 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_614
timestamp 1704896540
transform 1 0 57500 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_617
timestamp 1704896540
transform 1 0 57776 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_629
timestamp 1704896540
transform 1 0 58880 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_641
timestamp 1704896540
transform 1 0 59984 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_653
timestamp 1704896540
transform 1 0 61088 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_665
timestamp 1704896540
transform 1 0 62192 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_671
timestamp 1704896540
transform 1 0 62744 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_673
timestamp 1704896540
transform 1 0 62928 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_685
timestamp 1704896540
transform 1 0 64032 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_697
timestamp 1704896540
transform 1 0 65136 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_709
timestamp 1704896540
transform 1 0 66240 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_721
timestamp 1704896540
transform 1 0 67344 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_727
timestamp 1704896540
transform 1 0 67896 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_729
timestamp 1704896540
transform 1 0 68080 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_741
timestamp 1704896540
transform 1 0 69184 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_753
timestamp 1704896540
transform 1 0 70288 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_765
timestamp 1704896540
transform 1 0 71392 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_777
timestamp 1704896540
transform 1 0 72496 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_783
timestamp 1704896540
transform 1 0 73048 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_785
timestamp 1704896540
transform 1 0 73232 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_797
timestamp 1704896540
transform 1 0 74336 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1704896540
transform 1 0 1288 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1704896540
transform 1 0 2392 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1704896540
transform 1 0 3496 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1704896540
transform 1 0 3680 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1704896540
transform 1 0 4784 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1704896540
transform 1 0 5888 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1704896540
transform 1 0 6992 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1704896540
transform 1 0 8096 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1704896540
transform 1 0 8648 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1704896540
transform 1 0 8832 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1704896540
transform 1 0 9936 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1704896540
transform 1 0 11040 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1704896540
transform 1 0 12144 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1704896540
transform 1 0 13248 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1704896540
transform 1 0 13800 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1704896540
transform 1 0 13984 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1704896540
transform 1 0 15088 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1704896540
transform 1 0 16192 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1704896540
transform 1 0 17296 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1704896540
transform 1 0 18400 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1704896540
transform 1 0 18952 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1704896540
transform 1 0 19136 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1704896540
transform 1 0 20240 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1704896540
transform 1 0 21344 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1704896540
transform 1 0 22448 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 1704896540
transform 1 0 23552 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1704896540
transform 1 0 24104 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_253
timestamp 1704896540
transform 1 0 24288 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_263
timestamp 1704896540
transform 1 0 25208 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_282
timestamp 1704896540
transform 1 0 26956 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_309
timestamp 1704896540
transform 1 0 29440 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_337
timestamp 1704896540
transform 1 0 32016 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_377
timestamp 1704896540
transform 1 0 35696 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_391
timestamp 1704896540
transform 1 0 36984 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_397
timestamp 1704896540
transform 1 0 37536 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_404
timestamp 1704896540
transform 1 0 38180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_416
timestamp 1704896540
transform 1 0 39284 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_421
timestamp 1704896540
transform 1 0 39744 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_431
timestamp 1704896540
transform 1 0 40664 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_437
timestamp 1704896540
transform 1 0 41216 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_446
timestamp 1704896540
transform 1 0 42044 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_464
timestamp 1704896540
transform 1 0 43700 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_477
timestamp 1704896540
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_486
timestamp 1704896540
transform 1 0 45724 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_498
timestamp 1704896540
transform 1 0 46828 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_517
timestamp 1704896540
transform 1 0 48576 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_529
timestamp 1704896540
transform 1 0 49680 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_533
timestamp 1704896540
transform 1 0 50048 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_553
timestamp 1704896540
transform 1 0 51888 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_565
timestamp 1704896540
transform 1 0 52992 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_577
timestamp 1704896540
transform 1 0 54096 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_585
timestamp 1704896540
transform 1 0 54832 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_589
timestamp 1704896540
transform 1 0 55200 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_601
timestamp 1704896540
transform 1 0 56304 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_613
timestamp 1704896540
transform 1 0 57408 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_625
timestamp 1704896540
transform 1 0 58512 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_637
timestamp 1704896540
transform 1 0 59616 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_643
timestamp 1704896540
transform 1 0 60168 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_645
timestamp 1704896540
transform 1 0 60352 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_657
timestamp 1704896540
transform 1 0 61456 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_669
timestamp 1704896540
transform 1 0 62560 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_681
timestamp 1704896540
transform 1 0 63664 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_693
timestamp 1704896540
transform 1 0 64768 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_699
timestamp 1704896540
transform 1 0 65320 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_701
timestamp 1704896540
transform 1 0 65504 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_713
timestamp 1704896540
transform 1 0 66608 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_725
timestamp 1704896540
transform 1 0 67712 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_737
timestamp 1704896540
transform 1 0 68816 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_749
timestamp 1704896540
transform 1 0 69920 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_755
timestamp 1704896540
transform 1 0 70472 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_757
timestamp 1704896540
transform 1 0 70656 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_769
timestamp 1704896540
transform 1 0 71760 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_781
timestamp 1704896540
transform 1 0 72864 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_793
timestamp 1704896540
transform 1 0 73968 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1704896540
transform 1 0 1288 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1704896540
transform 1 0 2392 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1704896540
transform 1 0 3496 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1704896540
transform 1 0 4600 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1704896540
transform 1 0 5704 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1704896540
transform 1 0 6072 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1704896540
transform 1 0 6256 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1704896540
transform 1 0 7360 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1704896540
transform 1 0 8464 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1704896540
transform 1 0 9568 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1704896540
transform 1 0 10672 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1704896540
transform 1 0 11224 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1704896540
transform 1 0 11408 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1704896540
transform 1 0 12512 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1704896540
transform 1 0 13616 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1704896540
transform 1 0 14720 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1704896540
transform 1 0 15824 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1704896540
transform 1 0 16376 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1704896540
transform 1 0 16560 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1704896540
transform 1 0 17664 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 1704896540
transform 1 0 18768 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 1704896540
transform 1 0 19872 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1704896540
transform 1 0 20976 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1704896540
transform 1 0 21528 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1704896540
transform 1 0 21712 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1704896540
transform 1 0 22816 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 1704896540
transform 1 0 23920 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_261
timestamp 1704896540
transform 1 0 25024 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_269
timestamp 1704896540
transform 1 0 25760 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_289
timestamp 1704896540
transform 1 0 27600 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_300
timestamp 1704896540
transform 1 0 28612 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_323
timestamp 1704896540
transform 1 0 30728 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_334
timestamp 1704896540
transform 1 0 31740 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_343
timestamp 1704896540
transform 1 0 32568 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_354
timestamp 1704896540
transform 1 0 33580 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_366
timestamp 1704896540
transform 1 0 34684 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_378
timestamp 1704896540
transform 1 0 35788 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_390
timestamp 1704896540
transform 1 0 36892 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_401
timestamp 1704896540
transform 1 0 37904 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_407
timestamp 1704896540
transform 1 0 38456 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_416
timestamp 1704896540
transform 1 0 39284 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_424
timestamp 1704896540
transform 1 0 40020 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_433
timestamp 1704896540
transform 1 0 40848 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_439
timestamp 1704896540
transform 1 0 41400 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_469
timestamp 1704896540
transform 1 0 44160 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_491
timestamp 1704896540
transform 1 0 46184 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_495
timestamp 1704896540
transform 1 0 46552 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_505
timestamp 1704896540
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_514
timestamp 1704896540
transform 1 0 48300 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_555
timestamp 1704896540
transform 1 0 52072 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_559
timestamp 1704896540
transform 1 0 52440 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_609
timestamp 1704896540
transform 1 0 57040 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_615
timestamp 1704896540
transform 1 0 57592 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_617
timestamp 1704896540
transform 1 0 57776 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_629
timestamp 1704896540
transform 1 0 58880 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_641
timestamp 1704896540
transform 1 0 59984 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_653
timestamp 1704896540
transform 1 0 61088 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_665
timestamp 1704896540
transform 1 0 62192 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_671
timestamp 1704896540
transform 1 0 62744 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_673
timestamp 1704896540
transform 1 0 62928 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_685
timestamp 1704896540
transform 1 0 64032 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_697
timestamp 1704896540
transform 1 0 65136 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_709
timestamp 1704896540
transform 1 0 66240 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_721
timestamp 1704896540
transform 1 0 67344 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_727
timestamp 1704896540
transform 1 0 67896 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_729
timestamp 1704896540
transform 1 0 68080 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_741
timestamp 1704896540
transform 1 0 69184 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_753
timestamp 1704896540
transform 1 0 70288 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_765
timestamp 1704896540
transform 1 0 71392 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_777
timestamp 1704896540
transform 1 0 72496 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_783
timestamp 1704896540
transform 1 0 73048 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_785
timestamp 1704896540
transform 1 0 73232 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_797
timestamp 1704896540
transform 1 0 74336 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1704896540
transform 1 0 1288 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1704896540
transform 1 0 2392 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1704896540
transform 1 0 3496 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1704896540
transform 1 0 3680 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1704896540
transform 1 0 4784 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_53
timestamp 1704896540
transform 1 0 5888 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_57
timestamp 1704896540
transform 1 0 6256 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_69
timestamp 1704896540
transform 1 0 7360 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_81
timestamp 1704896540
transform 1 0 8464 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1704896540
transform 1 0 8832 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1704896540
transform 1 0 9936 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_109
timestamp 1704896540
transform 1 0 11040 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_113
timestamp 1704896540
transform 1 0 11408 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_125
timestamp 1704896540
transform 1 0 12512 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_137
timestamp 1704896540
transform 1 0 13616 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1704896540
transform 1 0 13984 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1704896540
transform 1 0 15088 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_165
timestamp 1704896540
transform 1 0 16192 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_169
timestamp 1704896540
transform 1 0 16560 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_181
timestamp 1704896540
transform 1 0 17664 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_193
timestamp 1704896540
transform 1 0 18768 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1704896540
transform 1 0 19136 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 1704896540
transform 1 0 20240 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_221
timestamp 1704896540
transform 1 0 21344 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_225
timestamp 1704896540
transform 1 0 21712 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_237
timestamp 1704896540
transform 1 0 22816 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_249
timestamp 1704896540
transform 1 0 23920 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1704896540
transform 1 0 24288 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 1704896540
transform 1 0 25392 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_277
timestamp 1704896540
transform 1 0 26496 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_281
timestamp 1704896540
transform 1 0 26864 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_293
timestamp 1704896540
transform 1 0 27968 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_301
timestamp 1704896540
transform 1 0 28704 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_323
timestamp 1704896540
transform 1 0 30728 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_332
timestamp 1704896540
transform 1 0 31556 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_337
timestamp 1704896540
transform 1 0 32016 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_349
timestamp 1704896540
transform 1 0 33120 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_361
timestamp 1704896540
transform 1 0 34224 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_365
timestamp 1704896540
transform 1 0 34592 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_391
timestamp 1704896540
transform 1 0 36984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_401
timestamp 1704896540
transform 1 0 37904 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_419
timestamp 1704896540
transform 1 0 39560 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_429
timestamp 1704896540
transform 1 0 40480 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_443
timestamp 1704896540
transform 1 0 41768 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_447
timestamp 1704896540
transform 1 0 42136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_473
timestamp 1704896540
transform 1 0 44528 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_477
timestamp 1704896540
transform 1 0 44896 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_483
timestamp 1704896540
transform 1 0 45448 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_500
timestamp 1704896540
transform 1 0 47012 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_529
timestamp 1704896540
transform 1 0 49680 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_557
timestamp 1704896540
transform 1 0 52256 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_561
timestamp 1704896540
transform 1 0 52624 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_573
timestamp 1704896540
transform 1 0 53728 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_579
timestamp 1704896540
transform 1 0 54280 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_613
timestamp 1704896540
transform 1 0 57408 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_617
timestamp 1704896540
transform 1 0 57776 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_629
timestamp 1704896540
transform 1 0 58880 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_633
timestamp 1704896540
transform 1 0 59248 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_642
timestamp 1704896540
transform 1 0 60076 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_653
timestamp 1704896540
transform 1 0 61088 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_665
timestamp 1704896540
transform 1 0 62192 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_671
timestamp 1704896540
transform 1 0 62744 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_673
timestamp 1704896540
transform 1 0 62928 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_685
timestamp 1704896540
transform 1 0 64032 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_697
timestamp 1704896540
transform 1 0 65136 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_701
timestamp 1704896540
transform 1 0 65504 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_713
timestamp 1704896540
transform 1 0 66608 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_725
timestamp 1704896540
transform 1 0 67712 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_729
timestamp 1704896540
transform 1 0 68080 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_741
timestamp 1704896540
transform 1 0 69184 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_753
timestamp 1704896540
transform 1 0 70288 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_757
timestamp 1704896540
transform 1 0 70656 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_769
timestamp 1704896540
transform 1 0 71760 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_781
timestamp 1704896540
transform 1 0 72864 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_785
timestamp 1704896540
transform 1 0 73232 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_797
timestamp 1704896540
transform 1 0 74336 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_702
timestamp 1704896540
transform 1 0 65596 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_714
timestamp 1704896540
transform 1 0 66700 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_726
timestamp 1704896540
transform 1 0 67804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_738
timestamp 1704896540
transform 1 0 68908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_750
timestamp 1704896540
transform 1 0 70012 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_754
timestamp 1704896540
transform 1 0 70380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_756
timestamp 1704896540
transform 1 0 70564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_768
timestamp 1704896540
transform 1 0 71668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_780
timestamp 1704896540
transform 1 0 72772 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_792
timestamp 1704896540
transform 1 0 73876 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_800
timestamp 1704896540
transform 1 0 74612 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_702
timestamp 1704896540
transform 1 0 65596 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_714
timestamp 1704896540
transform 1 0 66700 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_726
timestamp 1704896540
transform 1 0 67804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_728
timestamp 1704896540
transform 1 0 67988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_740
timestamp 1704896540
transform 1 0 69092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_752
timestamp 1704896540
transform 1 0 70196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_764
timestamp 1704896540
transform 1 0 71300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_776
timestamp 1704896540
transform 1 0 72404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_782
timestamp 1704896540
transform 1 0 72956 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_784
timestamp 1704896540
transform 1 0 73140 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_796
timestamp 1704896540
transform 1 0 74244 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_800
timestamp 1704896540
transform 1 0 74612 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_702
timestamp 1704896540
transform 1 0 65596 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_714
timestamp 1704896540
transform 1 0 66700 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_726
timestamp 1704896540
transform 1 0 67804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_738
timestamp 1704896540
transform 1 0 68908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_750
timestamp 1704896540
transform 1 0 70012 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_754
timestamp 1704896540
transform 1 0 70380 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_756
timestamp 1704896540
transform 1 0 70564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_768
timestamp 1704896540
transform 1 0 71668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_780
timestamp 1704896540
transform 1 0 72772 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_792
timestamp 1704896540
transform 1 0 73876 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_800
timestamp 1704896540
transform 1 0 74612 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_702
timestamp 1704896540
transform 1 0 65596 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_714
timestamp 1704896540
transform 1 0 66700 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_726
timestamp 1704896540
transform 1 0 67804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_728
timestamp 1704896540
transform 1 0 67988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_740
timestamp 1704896540
transform 1 0 69092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_752
timestamp 1704896540
transform 1 0 70196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_764
timestamp 1704896540
transform 1 0 71300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_776
timestamp 1704896540
transform 1 0 72404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_782
timestamp 1704896540
transform 1 0 72956 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_784
timestamp 1704896540
transform 1 0 73140 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_796
timestamp 1704896540
transform 1 0 74244 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_800
timestamp 1704896540
transform 1 0 74612 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_702
timestamp 1704896540
transform 1 0 65596 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_714
timestamp 1704896540
transform 1 0 66700 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_726
timestamp 1704896540
transform 1 0 67804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_738
timestamp 1704896540
transform 1 0 68908 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_750
timestamp 1704896540
transform 1 0 70012 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_754
timestamp 1704896540
transform 1 0 70380 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_756
timestamp 1704896540
transform 1 0 70564 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_768
timestamp 1704896540
transform 1 0 71668 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_780
timestamp 1704896540
transform 1 0 72772 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_792
timestamp 1704896540
transform 1 0 73876 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_800
timestamp 1704896540
transform 1 0 74612 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_702
timestamp 1704896540
transform 1 0 65596 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_714
timestamp 1704896540
transform 1 0 66700 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_726
timestamp 1704896540
transform 1 0 67804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_728
timestamp 1704896540
transform 1 0 67988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_740
timestamp 1704896540
transform 1 0 69092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_752
timestamp 1704896540
transform 1 0 70196 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_764
timestamp 1704896540
transform 1 0 71300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_776
timestamp 1704896540
transform 1 0 72404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_782
timestamp 1704896540
transform 1 0 72956 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_784
timestamp 1704896540
transform 1 0 73140 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_796
timestamp 1704896540
transform 1 0 74244 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_800
timestamp 1704896540
transform 1 0 74612 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_702
timestamp 1704896540
transform 1 0 65596 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_714
timestamp 1704896540
transform 1 0 66700 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_726
timestamp 1704896540
transform 1 0 67804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_738
timestamp 1704896540
transform 1 0 68908 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_750
timestamp 1704896540
transform 1 0 70012 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_754
timestamp 1704896540
transform 1 0 70380 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_756
timestamp 1704896540
transform 1 0 70564 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_768
timestamp 1704896540
transform 1 0 71668 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_780
timestamp 1704896540
transform 1 0 72772 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_792
timestamp 1704896540
transform 1 0 73876 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_800
timestamp 1704896540
transform 1 0 74612 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_702
timestamp 1704896540
transform 1 0 65596 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_714
timestamp 1704896540
transform 1 0 66700 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_726
timestamp 1704896540
transform 1 0 67804 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_728
timestamp 1704896540
transform 1 0 67988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_740
timestamp 1704896540
transform 1 0 69092 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_752
timestamp 1704896540
transform 1 0 70196 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_764
timestamp 1704896540
transform 1 0 71300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_776
timestamp 1704896540
transform 1 0 72404 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_782
timestamp 1704896540
transform 1 0 72956 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_784
timestamp 1704896540
transform 1 0 73140 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_796
timestamp 1704896540
transform 1 0 74244 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_800
timestamp 1704896540
transform 1 0 74612 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_702
timestamp 1704896540
transform 1 0 65596 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_714
timestamp 1704896540
transform 1 0 66700 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_726
timestamp 1704896540
transform 1 0 67804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_738
timestamp 1704896540
transform 1 0 68908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_750
timestamp 1704896540
transform 1 0 70012 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_754
timestamp 1704896540
transform 1 0 70380 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_756
timestamp 1704896540
transform 1 0 70564 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_768
timestamp 1704896540
transform 1 0 71668 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_780
timestamp 1704896540
transform 1 0 72772 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_792
timestamp 1704896540
transform 1 0 73876 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_800
timestamp 1704896540
transform 1 0 74612 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_702
timestamp 1704896540
transform 1 0 65596 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_714
timestamp 1704896540
transform 1 0 66700 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_726
timestamp 1704896540
transform 1 0 67804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_728
timestamp 1704896540
transform 1 0 67988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_740
timestamp 1704896540
transform 1 0 69092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_752
timestamp 1704896540
transform 1 0 70196 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_764
timestamp 1704896540
transform 1 0 71300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_776
timestamp 1704896540
transform 1 0 72404 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_782
timestamp 1704896540
transform 1 0 72956 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_784
timestamp 1704896540
transform 1 0 73140 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_796
timestamp 1704896540
transform 1 0 74244 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_800
timestamp 1704896540
transform 1 0 74612 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_710
timestamp 1704896540
transform 1 0 66332 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_722
timestamp 1704896540
transform 1 0 67436 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_734
timestamp 1704896540
transform 1 0 68540 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_746
timestamp 1704896540
transform 1 0 69644 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_754
timestamp 1704896540
transform 1 0 70380 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_756
timestamp 1704896540
transform 1 0 70564 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_768
timestamp 1704896540
transform 1 0 71668 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_780
timestamp 1704896540
transform 1 0 72772 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_792
timestamp 1704896540
transform 1 0 73876 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_800
timestamp 1704896540
transform 1 0 74612 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_702
timestamp 1704896540
transform 1 0 65596 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_714
timestamp 1704896540
transform 1 0 66700 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_726
timestamp 1704896540
transform 1 0 67804 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_728
timestamp 1704896540
transform 1 0 67988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_740
timestamp 1704896540
transform 1 0 69092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_752
timestamp 1704896540
transform 1 0 70196 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_764
timestamp 1704896540
transform 1 0 71300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_776
timestamp 1704896540
transform 1 0 72404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_782
timestamp 1704896540
transform 1 0 72956 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_784
timestamp 1704896540
transform 1 0 73140 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_796
timestamp 1704896540
transform 1 0 74244 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_800
timestamp 1704896540
transform 1 0 74612 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_702
timestamp 1704896540
transform 1 0 65596 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_714
timestamp 1704896540
transform 1 0 66700 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_726
timestamp 1704896540
transform 1 0 67804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_738
timestamp 1704896540
transform 1 0 68908 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_750
timestamp 1704896540
transform 1 0 70012 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_754
timestamp 1704896540
transform 1 0 70380 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_756
timestamp 1704896540
transform 1 0 70564 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_768
timestamp 1704896540
transform 1 0 71668 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_780
timestamp 1704896540
transform 1 0 72772 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_792
timestamp 1704896540
transform 1 0 73876 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_800
timestamp 1704896540
transform 1 0 74612 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_710
timestamp 1704896540
transform 1 0 66332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_722
timestamp 1704896540
transform 1 0 67436 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_726
timestamp 1704896540
transform 1 0 67804 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_728
timestamp 1704896540
transform 1 0 67988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_740
timestamp 1704896540
transform 1 0 69092 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_752
timestamp 1704896540
transform 1 0 70196 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_764
timestamp 1704896540
transform 1 0 71300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_776
timestamp 1704896540
transform 1 0 72404 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_782
timestamp 1704896540
transform 1 0 72956 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_784
timestamp 1704896540
transform 1 0 73140 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_796
timestamp 1704896540
transform 1 0 74244 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_800
timestamp 1704896540
transform 1 0 74612 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_702
timestamp 1704896540
transform 1 0 65596 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_714
timestamp 1704896540
transform 1 0 66700 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_726
timestamp 1704896540
transform 1 0 67804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_738
timestamp 1704896540
transform 1 0 68908 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_750
timestamp 1704896540
transform 1 0 70012 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_754
timestamp 1704896540
transform 1 0 70380 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_756
timestamp 1704896540
transform 1 0 70564 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_768
timestamp 1704896540
transform 1 0 71668 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_780
timestamp 1704896540
transform 1 0 72772 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_792
timestamp 1704896540
transform 1 0 73876 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_800
timestamp 1704896540
transform 1 0 74612 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_710
timestamp 1704896540
transform 1 0 66332 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_722
timestamp 1704896540
transform 1 0 67436 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_726
timestamp 1704896540
transform 1 0 67804 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_728
timestamp 1704896540
transform 1 0 67988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_740
timestamp 1704896540
transform 1 0 69092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_752
timestamp 1704896540
transform 1 0 70196 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_764
timestamp 1704896540
transform 1 0 71300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_776
timestamp 1704896540
transform 1 0 72404 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_782
timestamp 1704896540
transform 1 0 72956 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_784
timestamp 1704896540
transform 1 0 73140 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_796
timestamp 1704896540
transform 1 0 74244 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_800
timestamp 1704896540
transform 1 0 74612 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_710
timestamp 1704896540
transform 1 0 66332 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_722
timestamp 1704896540
transform 1 0 67436 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_734
timestamp 1704896540
transform 1 0 68540 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_746
timestamp 1704896540
transform 1 0 69644 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_754
timestamp 1704896540
transform 1 0 70380 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_756
timestamp 1704896540
transform 1 0 70564 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_768
timestamp 1704896540
transform 1 0 71668 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_780
timestamp 1704896540
transform 1 0 72772 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_792
timestamp 1704896540
transform 1 0 73876 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_800
timestamp 1704896540
transform 1 0 74612 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_710
timestamp 1704896540
transform 1 0 66332 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_722
timestamp 1704896540
transform 1 0 67436 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_726
timestamp 1704896540
transform 1 0 67804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_728
timestamp 1704896540
transform 1 0 67988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_740
timestamp 1704896540
transform 1 0 69092 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_752
timestamp 1704896540
transform 1 0 70196 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_764
timestamp 1704896540
transform 1 0 71300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_776
timestamp 1704896540
transform 1 0 72404 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_782
timestamp 1704896540
transform 1 0 72956 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_784
timestamp 1704896540
transform 1 0 73140 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_796
timestamp 1704896540
transform 1 0 74244 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_800
timestamp 1704896540
transform 1 0 74612 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_710
timestamp 1704896540
transform 1 0 66332 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_722
timestamp 1704896540
transform 1 0 67436 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_734
timestamp 1704896540
transform 1 0 68540 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_746
timestamp 1704896540
transform 1 0 69644 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_754
timestamp 1704896540
transform 1 0 70380 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_756
timestamp 1704896540
transform 1 0 70564 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_768
timestamp 1704896540
transform 1 0 71668 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_780
timestamp 1704896540
transform 1 0 72772 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_792
timestamp 1704896540
transform 1 0 73876 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_800
timestamp 1704896540
transform 1 0 74612 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_710
timestamp 1704896540
transform 1 0 66332 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_722
timestamp 1704896540
transform 1 0 67436 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_726
timestamp 1704896540
transform 1 0 67804 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_728
timestamp 1704896540
transform 1 0 67988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_740
timestamp 1704896540
transform 1 0 69092 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_752
timestamp 1704896540
transform 1 0 70196 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_764
timestamp 1704896540
transform 1 0 71300 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_776
timestamp 1704896540
transform 1 0 72404 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_782
timestamp 1704896540
transform 1 0 72956 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_784
timestamp 1704896540
transform 1 0 73140 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_796
timestamp 1704896540
transform 1 0 74244 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_800
timestamp 1704896540
transform 1 0 74612 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_718
timestamp 1704896540
transform 1 0 67068 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_730
timestamp 1704896540
transform 1 0 68172 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_742
timestamp 1704896540
transform 1 0 69276 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_754
timestamp 1704896540
transform 1 0 70380 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_756
timestamp 1704896540
transform 1 0 70564 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_768
timestamp 1704896540
transform 1 0 71668 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_780
timestamp 1704896540
transform 1 0 72772 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_792
timestamp 1704896540
transform 1 0 73876 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_800
timestamp 1704896540
transform 1 0 74612 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_710
timestamp 1704896540
transform 1 0 66332 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_722
timestamp 1704896540
transform 1 0 67436 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_726
timestamp 1704896540
transform 1 0 67804 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_728
timestamp 1704896540
transform 1 0 67988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_740
timestamp 1704896540
transform 1 0 69092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_752
timestamp 1704896540
transform 1 0 70196 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_764
timestamp 1704896540
transform 1 0 71300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_776
timestamp 1704896540
transform 1 0 72404 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_782
timestamp 1704896540
transform 1 0 72956 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_784
timestamp 1704896540
transform 1 0 73140 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_796
timestamp 1704896540
transform 1 0 74244 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_800
timestamp 1704896540
transform 1 0 74612 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_710
timestamp 1704896540
transform 1 0 66332 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_722
timestamp 1704896540
transform 1 0 67436 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_734
timestamp 1704896540
transform 1 0 68540 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_746
timestamp 1704896540
transform 1 0 69644 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_754
timestamp 1704896540
transform 1 0 70380 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_756
timestamp 1704896540
transform 1 0 70564 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_768
timestamp 1704896540
transform 1 0 71668 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_780
timestamp 1704896540
transform 1 0 72772 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_792
timestamp 1704896540
transform 1 0 73876 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_800
timestamp 1704896540
transform 1 0 74612 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_710
timestamp 1704896540
transform 1 0 66332 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_722
timestamp 1704896540
transform 1 0 67436 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_726
timestamp 1704896540
transform 1 0 67804 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_728
timestamp 1704896540
transform 1 0 67988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_740
timestamp 1704896540
transform 1 0 69092 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_752
timestamp 1704896540
transform 1 0 70196 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_764
timestamp 1704896540
transform 1 0 71300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_776
timestamp 1704896540
transform 1 0 72404 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_782
timestamp 1704896540
transform 1 0 72956 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_784
timestamp 1704896540
transform 1 0 73140 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_796
timestamp 1704896540
transform 1 0 74244 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_800
timestamp 1704896540
transform 1 0 74612 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_710
timestamp 1704896540
transform 1 0 66332 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_722
timestamp 1704896540
transform 1 0 67436 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_734
timestamp 1704896540
transform 1 0 68540 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_746
timestamp 1704896540
transform 1 0 69644 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_754
timestamp 1704896540
transform 1 0 70380 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_756
timestamp 1704896540
transform 1 0 70564 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_768
timestamp 1704896540
transform 1 0 71668 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_780
timestamp 1704896540
transform 1 0 72772 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_792
timestamp 1704896540
transform 1 0 73876 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_800
timestamp 1704896540
transform 1 0 74612 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_710
timestamp 1704896540
transform 1 0 66332 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_722
timestamp 1704896540
transform 1 0 67436 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_726
timestamp 1704896540
transform 1 0 67804 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_728
timestamp 1704896540
transform 1 0 67988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_740
timestamp 1704896540
transform 1 0 69092 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_752
timestamp 1704896540
transform 1 0 70196 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_764
timestamp 1704896540
transform 1 0 71300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_776
timestamp 1704896540
transform 1 0 72404 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_782
timestamp 1704896540
transform 1 0 72956 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_784
timestamp 1704896540
transform 1 0 73140 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_796
timestamp 1704896540
transform 1 0 74244 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_800
timestamp 1704896540
transform 1 0 74612 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_726
timestamp 1704896540
transform 1 0 67804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_738
timestamp 1704896540
transform 1 0 68908 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_750
timestamp 1704896540
transform 1 0 70012 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_754
timestamp 1704896540
transform 1 0 70380 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_756
timestamp 1704896540
transform 1 0 70564 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_768
timestamp 1704896540
transform 1 0 71668 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_780
timestamp 1704896540
transform 1 0 72772 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_792
timestamp 1704896540
transform 1 0 73876 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_800
timestamp 1704896540
transform 1 0 74612 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_702
timestamp 1704896540
transform 1 0 65596 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_714
timestamp 1704896540
transform 1 0 66700 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_726
timestamp 1704896540
transform 1 0 67804 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_728
timestamp 1704896540
transform 1 0 67988 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_738
timestamp 1704896540
transform 1 0 68908 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_750
timestamp 1704896540
transform 1 0 70012 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_762
timestamp 1704896540
transform 1 0 71116 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_774
timestamp 1704896540
transform 1 0 72220 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_782
timestamp 1704896540
transform 1 0 72956 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_784
timestamp 1704896540
transform 1 0 73140 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_796
timestamp 1704896540
transform 1 0 74244 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_800
timestamp 1704896540
transform 1 0 74612 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_710
timestamp 1704896540
transform 1 0 66332 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_722
timestamp 1704896540
transform 1 0 67436 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_734
timestamp 1704896540
transform 1 0 68540 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_746
timestamp 1704896540
transform 1 0 69644 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_754
timestamp 1704896540
transform 1 0 70380 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_756
timestamp 1704896540
transform 1 0 70564 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_768
timestamp 1704896540
transform 1 0 71668 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_780
timestamp 1704896540
transform 1 0 72772 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_792
timestamp 1704896540
transform 1 0 73876 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_800
timestamp 1704896540
transform 1 0 74612 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_718
timestamp 1704896540
transform 1 0 67068 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_726
timestamp 1704896540
transform 1 0 67804 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_728
timestamp 1704896540
transform 1 0 67988 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_734
timestamp 1704896540
transform 1 0 68540 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_743
timestamp 1704896540
transform 1 0 69368 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_759
timestamp 1704896540
transform 1 0 70840 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_771
timestamp 1704896540
transform 1 0 71944 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_784
timestamp 1704896540
transform 1 0 73140 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_796
timestamp 1704896540
transform 1 0 74244 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_800
timestamp 1704896540
transform 1 0 74612 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_710
timestamp 1704896540
transform 1 0 66332 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_722
timestamp 1704896540
transform 1 0 67436 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_734
timestamp 1704896540
transform 1 0 68540 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_746
timestamp 1704896540
transform 1 0 69644 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_754
timestamp 1704896540
transform 1 0 70380 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_756
timestamp 1704896540
transform 1 0 70564 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_768
timestamp 1704896540
transform 1 0 71668 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_780
timestamp 1704896540
transform 1 0 72772 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_792
timestamp 1704896540
transform 1 0 73876 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_800
timestamp 1704896540
transform 1 0 74612 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_726
timestamp 1704896540
transform 1 0 67804 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_728
timestamp 1704896540
transform 1 0 67988 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_740
timestamp 1704896540
transform 1 0 69092 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_752
timestamp 1704896540
transform 1 0 70196 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_764
timestamp 1704896540
transform 1 0 71300 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_776
timestamp 1704896540
transform 1 0 72404 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_782
timestamp 1704896540
transform 1 0 72956 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_784
timestamp 1704896540
transform 1 0 73140 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_796
timestamp 1704896540
transform 1 0 74244 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_800
timestamp 1704896540
transform 1 0 74612 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_726
timestamp 1704896540
transform 1 0 67804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_738
timestamp 1704896540
transform 1 0 68908 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_750
timestamp 1704896540
transform 1 0 70012 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_754
timestamp 1704896540
transform 1 0 70380 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_756
timestamp 1704896540
transform 1 0 70564 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_768
timestamp 1704896540
transform 1 0 71668 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_780
timestamp 1704896540
transform 1 0 72772 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_792
timestamp 1704896540
transform 1 0 73876 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_800
timestamp 1704896540
transform 1 0 74612 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_718
timestamp 1704896540
transform 1 0 67068 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_726
timestamp 1704896540
transform 1 0 67804 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_728
timestamp 1704896540
transform 1 0 67988 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_740
timestamp 1704896540
transform 1 0 69092 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_752
timestamp 1704896540
transform 1 0 70196 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_764
timestamp 1704896540
transform 1 0 71300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_776
timestamp 1704896540
transform 1 0 72404 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_782
timestamp 1704896540
transform 1 0 72956 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_784
timestamp 1704896540
transform 1 0 73140 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_796
timestamp 1704896540
transform 1 0 74244 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_800
timestamp 1704896540
transform 1 0 74612 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_718
timestamp 1704896540
transform 1 0 67068 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_730
timestamp 1704896540
transform 1 0 68172 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_742
timestamp 1704896540
transform 1 0 69276 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_754
timestamp 1704896540
transform 1 0 70380 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_756
timestamp 1704896540
transform 1 0 70564 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_768
timestamp 1704896540
transform 1 0 71668 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_780
timestamp 1704896540
transform 1 0 72772 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_792
timestamp 1704896540
transform 1 0 73876 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_800
timestamp 1704896540
transform 1 0 74612 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_710
timestamp 1704896540
transform 1 0 66332 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_722
timestamp 1704896540
transform 1 0 67436 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_726
timestamp 1704896540
transform 1 0 67804 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_728
timestamp 1704896540
transform 1 0 67988 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_740
timestamp 1704896540
transform 1 0 69092 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_752
timestamp 1704896540
transform 1 0 70196 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_764
timestamp 1704896540
transform 1 0 71300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_776
timestamp 1704896540
transform 1 0 72404 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_782
timestamp 1704896540
transform 1 0 72956 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_784
timestamp 1704896540
transform 1 0 73140 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_796
timestamp 1704896540
transform 1 0 74244 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_800
timestamp 1704896540
transform 1 0 74612 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_710
timestamp 1704896540
transform 1 0 66332 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_722
timestamp 1704896540
transform 1 0 67436 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_734
timestamp 1704896540
transform 1 0 68540 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_746
timestamp 1704896540
transform 1 0 69644 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_754
timestamp 1704896540
transform 1 0 70380 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_756
timestamp 1704896540
transform 1 0 70564 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_768
timestamp 1704896540
transform 1 0 71668 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_780
timestamp 1704896540
transform 1 0 72772 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_792
timestamp 1704896540
transform 1 0 73876 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_800
timestamp 1704896540
transform 1 0 74612 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_710
timestamp 1704896540
transform 1 0 66332 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_722
timestamp 1704896540
transform 1 0 67436 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_726
timestamp 1704896540
transform 1 0 67804 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_728
timestamp 1704896540
transform 1 0 67988 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_740
timestamp 1704896540
transform 1 0 69092 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_752
timestamp 1704896540
transform 1 0 70196 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_764
timestamp 1704896540
transform 1 0 71300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_776
timestamp 1704896540
transform 1 0 72404 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_782
timestamp 1704896540
transform 1 0 72956 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_784
timestamp 1704896540
transform 1 0 73140 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_796
timestamp 1704896540
transform 1 0 74244 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_800
timestamp 1704896540
transform 1 0 74612 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_726
timestamp 1704896540
transform 1 0 67804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_738
timestamp 1704896540
transform 1 0 68908 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_750
timestamp 1704896540
transform 1 0 70012 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_754
timestamp 1704896540
transform 1 0 70380 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_756
timestamp 1704896540
transform 1 0 70564 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_768
timestamp 1704896540
transform 1 0 71668 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_780
timestamp 1704896540
transform 1 0 72772 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_792
timestamp 1704896540
transform 1 0 73876 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_800
timestamp 1704896540
transform 1 0 74612 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_718
timestamp 1704896540
transform 1 0 67068 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_726
timestamp 1704896540
transform 1 0 67804 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_728
timestamp 1704896540
transform 1 0 67988 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_740
timestamp 1704896540
transform 1 0 69092 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_752
timestamp 1704896540
transform 1 0 70196 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_764
timestamp 1704896540
transform 1 0 71300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_776
timestamp 1704896540
transform 1 0 72404 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_782
timestamp 1704896540
transform 1 0 72956 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_784
timestamp 1704896540
transform 1 0 73140 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_796
timestamp 1704896540
transform 1 0 74244 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_800
timestamp 1704896540
transform 1 0 74612 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_710
timestamp 1704896540
transform 1 0 66332 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_714
timestamp 1704896540
transform 1 0 66700 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_726
timestamp 1704896540
transform 1 0 67804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_738
timestamp 1704896540
transform 1 0 68908 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_750
timestamp 1704896540
transform 1 0 70012 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_754
timestamp 1704896540
transform 1 0 70380 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_756
timestamp 1704896540
transform 1 0 70564 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_768
timestamp 1704896540
transform 1 0 71668 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_780
timestamp 1704896540
transform 1 0 72772 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_792
timestamp 1704896540
transform 1 0 73876 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_800
timestamp 1704896540
transform 1 0 74612 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_722
timestamp 1704896540
transform 1 0 67436 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_726
timestamp 1704896540
transform 1 0 67804 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_728
timestamp 1704896540
transform 1 0 67988 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_740
timestamp 1704896540
transform 1 0 69092 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_752
timestamp 1704896540
transform 1 0 70196 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_764
timestamp 1704896540
transform 1 0 71300 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_776
timestamp 1704896540
transform 1 0 72404 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_782
timestamp 1704896540
transform 1 0 72956 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_784
timestamp 1704896540
transform 1 0 73140 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_796
timestamp 1704896540
transform 1 0 74244 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_800
timestamp 1704896540
transform 1 0 74612 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_710
timestamp 1704896540
transform 1 0 66332 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_722
timestamp 1704896540
transform 1 0 67436 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_734
timestamp 1704896540
transform 1 0 68540 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_746
timestamp 1704896540
transform 1 0 69644 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_754
timestamp 1704896540
transform 1 0 70380 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_756
timestamp 1704896540
transform 1 0 70564 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_768
timestamp 1704896540
transform 1 0 71668 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_780
timestamp 1704896540
transform 1 0 72772 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_792
timestamp 1704896540
transform 1 0 73876 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_800
timestamp 1704896540
transform 1 0 74612 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_710
timestamp 1704896540
transform 1 0 66332 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_722
timestamp 1704896540
transform 1 0 67436 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_726
timestamp 1704896540
transform 1 0 67804 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_728
timestamp 1704896540
transform 1 0 67988 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_740
timestamp 1704896540
transform 1 0 69092 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_752
timestamp 1704896540
transform 1 0 70196 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_764
timestamp 1704896540
transform 1 0 71300 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_776
timestamp 1704896540
transform 1 0 72404 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_782
timestamp 1704896540
transform 1 0 72956 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_784
timestamp 1704896540
transform 1 0 73140 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_796
timestamp 1704896540
transform 1 0 74244 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_800
timestamp 1704896540
transform 1 0 74612 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_710
timestamp 1704896540
transform 1 0 66332 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_722
timestamp 1704896540
transform 1 0 67436 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_734
timestamp 1704896540
transform 1 0 68540 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_746
timestamp 1704896540
transform 1 0 69644 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_754
timestamp 1704896540
transform 1 0 70380 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_756
timestamp 1704896540
transform 1 0 70564 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_768
timestamp 1704896540
transform 1 0 71668 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_780
timestamp 1704896540
transform 1 0 72772 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_792
timestamp 1704896540
transform 1 0 73876 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_800
timestamp 1704896540
transform 1 0 74612 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_710
timestamp 1704896540
transform 1 0 66332 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_722
timestamp 1704896540
transform 1 0 67436 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_726
timestamp 1704896540
transform 1 0 67804 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_728
timestamp 1704896540
transform 1 0 67988 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_740
timestamp 1704896540
transform 1 0 69092 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_752
timestamp 1704896540
transform 1 0 70196 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_764
timestamp 1704896540
transform 1 0 71300 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_776
timestamp 1704896540
transform 1 0 72404 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_782
timestamp 1704896540
transform 1 0 72956 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_784
timestamp 1704896540
transform 1 0 73140 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_796
timestamp 1704896540
transform 1 0 74244 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_800
timestamp 1704896540
transform 1 0 74612 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_710
timestamp 1704896540
transform 1 0 66332 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_722
timestamp 1704896540
transform 1 0 67436 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_734
timestamp 1704896540
transform 1 0 68540 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_746
timestamp 1704896540
transform 1 0 69644 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_754
timestamp 1704896540
transform 1 0 70380 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_756
timestamp 1704896540
transform 1 0 70564 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_768
timestamp 1704896540
transform 1 0 71668 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_780
timestamp 1704896540
transform 1 0 72772 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_792
timestamp 1704896540
transform 1 0 73876 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_800
timestamp 1704896540
transform 1 0 74612 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_710
timestamp 1704896540
transform 1 0 66332 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_722
timestamp 1704896540
transform 1 0 67436 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_726
timestamp 1704896540
transform 1 0 67804 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_728
timestamp 1704896540
transform 1 0 67988 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_740
timestamp 1704896540
transform 1 0 69092 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_752
timestamp 1704896540
transform 1 0 70196 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_764
timestamp 1704896540
transform 1 0 71300 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_776
timestamp 1704896540
transform 1 0 72404 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_782
timestamp 1704896540
transform 1 0 72956 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_784
timestamp 1704896540
transform 1 0 73140 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_796
timestamp 1704896540
transform 1 0 74244 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_800
timestamp 1704896540
transform 1 0 74612 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_710
timestamp 1704896540
transform 1 0 66332 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_722
timestamp 1704896540
transform 1 0 67436 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_734
timestamp 1704896540
transform 1 0 68540 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_746
timestamp 1704896540
transform 1 0 69644 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_754
timestamp 1704896540
transform 1 0 70380 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_756
timestamp 1704896540
transform 1 0 70564 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_768
timestamp 1704896540
transform 1 0 71668 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_780
timestamp 1704896540
transform 1 0 72772 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_792
timestamp 1704896540
transform 1 0 73876 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_800
timestamp 1704896540
transform 1 0 74612 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_710
timestamp 1704896540
transform 1 0 66332 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_722
timestamp 1704896540
transform 1 0 67436 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_726
timestamp 1704896540
transform 1 0 67804 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_728
timestamp 1704896540
transform 1 0 67988 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_740
timestamp 1704896540
transform 1 0 69092 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_752
timestamp 1704896540
transform 1 0 70196 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_764
timestamp 1704896540
transform 1 0 71300 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_776
timestamp 1704896540
transform 1 0 72404 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_782
timestamp 1704896540
transform 1 0 72956 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_784
timestamp 1704896540
transform 1 0 73140 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_796
timestamp 1704896540
transform 1 0 74244 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_800
timestamp 1704896540
transform 1 0 74612 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_710
timestamp 1704896540
transform 1 0 66332 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_722
timestamp 1704896540
transform 1 0 67436 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_734
timestamp 1704896540
transform 1 0 68540 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_746
timestamp 1704896540
transform 1 0 69644 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_754
timestamp 1704896540
transform 1 0 70380 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_756
timestamp 1704896540
transform 1 0 70564 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_768
timestamp 1704896540
transform 1 0 71668 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_780
timestamp 1704896540
transform 1 0 72772 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_792
timestamp 1704896540
transform 1 0 73876 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_800
timestamp 1704896540
transform 1 0 74612 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_726
timestamp 1704896540
transform 1 0 67804 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_728
timestamp 1704896540
transform 1 0 67988 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_740
timestamp 1704896540
transform 1 0 69092 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_752
timestamp 1704896540
transform 1 0 70196 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_764
timestamp 1704896540
transform 1 0 71300 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_776
timestamp 1704896540
transform 1 0 72404 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_782
timestamp 1704896540
transform 1 0 72956 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_784
timestamp 1704896540
transform 1 0 73140 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_796
timestamp 1704896540
transform 1 0 74244 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_800
timestamp 1704896540
transform 1 0 74612 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_726
timestamp 1704896540
transform 1 0 67804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_738
timestamp 1704896540
transform 1 0 68908 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_750
timestamp 1704896540
transform 1 0 70012 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_754
timestamp 1704896540
transform 1 0 70380 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_756
timestamp 1704896540
transform 1 0 70564 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_768
timestamp 1704896540
transform 1 0 71668 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_780
timestamp 1704896540
transform 1 0 72772 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_792
timestamp 1704896540
transform 1 0 73876 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_800
timestamp 1704896540
transform 1 0 74612 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_722
timestamp 1704896540
transform 1 0 67436 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_726
timestamp 1704896540
transform 1 0 67804 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_736
timestamp 1704896540
transform 1 0 68724 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_748
timestamp 1704896540
transform 1 0 69828 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_760
timestamp 1704896540
transform 1 0 70932 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_772
timestamp 1704896540
transform 1 0 72036 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_780
timestamp 1704896540
transform 1 0 72772 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_784
timestamp 1704896540
transform 1 0 73140 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_796
timestamp 1704896540
transform 1 0 74244 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_800
timestamp 1704896540
transform 1 0 74612 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_726
timestamp 1704896540
transform 1 0 67804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_738
timestamp 1704896540
transform 1 0 68908 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_750
timestamp 1704896540
transform 1 0 70012 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_754
timestamp 1704896540
transform 1 0 70380 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_756
timestamp 1704896540
transform 1 0 70564 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_768
timestamp 1704896540
transform 1 0 71668 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_780
timestamp 1704896540
transform 1 0 72772 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_792
timestamp 1704896540
transform 1 0 73876 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_800
timestamp 1704896540
transform 1 0 74612 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_718
timestamp 1704896540
transform 1 0 67068 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_726
timestamp 1704896540
transform 1 0 67804 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_728
timestamp 1704896540
transform 1 0 67988 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_740
timestamp 1704896540
transform 1 0 69092 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_752
timestamp 1704896540
transform 1 0 70196 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_764
timestamp 1704896540
transform 1 0 71300 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_776
timestamp 1704896540
transform 1 0 72404 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_782
timestamp 1704896540
transform 1 0 72956 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_784
timestamp 1704896540
transform 1 0 73140 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_796
timestamp 1704896540
transform 1 0 74244 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_800
timestamp 1704896540
transform 1 0 74612 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_710
timestamp 1704896540
transform 1 0 66332 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_722
timestamp 1704896540
transform 1 0 67436 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_734
timestamp 1704896540
transform 1 0 68540 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_746
timestamp 1704896540
transform 1 0 69644 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_754
timestamp 1704896540
transform 1 0 70380 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_756
timestamp 1704896540
transform 1 0 70564 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_768
timestamp 1704896540
transform 1 0 71668 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_780
timestamp 1704896540
transform 1 0 72772 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_792
timestamp 1704896540
transform 1 0 73876 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_800
timestamp 1704896540
transform 1 0 74612 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_710
timestamp 1704896540
transform 1 0 66332 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_722
timestamp 1704896540
transform 1 0 67436 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_726
timestamp 1704896540
transform 1 0 67804 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_728
timestamp 1704896540
transform 1 0 67988 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_740
timestamp 1704896540
transform 1 0 69092 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_752
timestamp 1704896540
transform 1 0 70196 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_764
timestamp 1704896540
transform 1 0 71300 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_776
timestamp 1704896540
transform 1 0 72404 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_782
timestamp 1704896540
transform 1 0 72956 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_784
timestamp 1704896540
transform 1 0 73140 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_796
timestamp 1704896540
transform 1 0 74244 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_800
timestamp 1704896540
transform 1 0 74612 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_710
timestamp 1704896540
transform 1 0 66332 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_722
timestamp 1704896540
transform 1 0 67436 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_734
timestamp 1704896540
transform 1 0 68540 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_746
timestamp 1704896540
transform 1 0 69644 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_754
timestamp 1704896540
transform 1 0 70380 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_756
timestamp 1704896540
transform 1 0 70564 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_768
timestamp 1704896540
transform 1 0 71668 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_780
timestamp 1704896540
transform 1 0 72772 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_792
timestamp 1704896540
transform 1 0 73876 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_800
timestamp 1704896540
transform 1 0 74612 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_710
timestamp 1704896540
transform 1 0 66332 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68_722
timestamp 1704896540
transform 1 0 67436 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_726
timestamp 1704896540
transform 1 0 67804 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_728
timestamp 1704896540
transform 1 0 67988 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_740
timestamp 1704896540
transform 1 0 69092 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_752
timestamp 1704896540
transform 1 0 70196 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_764
timestamp 1704896540
transform 1 0 71300 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_776
timestamp 1704896540
transform 1 0 72404 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_782
timestamp 1704896540
transform 1 0 72956 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_784
timestamp 1704896540
transform 1 0 73140 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68_796
timestamp 1704896540
transform 1 0 74244 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_800
timestamp 1704896540
transform 1 0 74612 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_710
timestamp 1704896540
transform 1 0 66332 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_722
timestamp 1704896540
transform 1 0 67436 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_734
timestamp 1704896540
transform 1 0 68540 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69_746
timestamp 1704896540
transform 1 0 69644 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_754
timestamp 1704896540
transform 1 0 70380 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_756
timestamp 1704896540
transform 1 0 70564 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_768
timestamp 1704896540
transform 1 0 71668 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_780
timestamp 1704896540
transform 1 0 72772 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69_792
timestamp 1704896540
transform 1 0 73876 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_800
timestamp 1704896540
transform 1 0 74612 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_710
timestamp 1704896540
transform 1 0 66332 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_70_722
timestamp 1704896540
transform 1 0 67436 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_726
timestamp 1704896540
transform 1 0 67804 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_728
timestamp 1704896540
transform 1 0 67988 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_740
timestamp 1704896540
transform 1 0 69092 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_752
timestamp 1704896540
transform 1 0 70196 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_764
timestamp 1704896540
transform 1 0 71300 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_776
timestamp 1704896540
transform 1 0 72404 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_782
timestamp 1704896540
transform 1 0 72956 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_784
timestamp 1704896540
transform 1 0 73140 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_70_796
timestamp 1704896540
transform 1 0 74244 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_800
timestamp 1704896540
transform 1 0 74612 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_710
timestamp 1704896540
transform 1 0 66332 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_722
timestamp 1704896540
transform 1 0 67436 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_734
timestamp 1704896540
transform 1 0 68540 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_71_746
timestamp 1704896540
transform 1 0 69644 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_754
timestamp 1704896540
transform 1 0 70380 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_756
timestamp 1704896540
transform 1 0 70564 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_768
timestamp 1704896540
transform 1 0 71668 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_780
timestamp 1704896540
transform 1 0 72772 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_71_792
timestamp 1704896540
transform 1 0 73876 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_800
timestamp 1704896540
transform 1 0 74612 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_726
timestamp 1704896540
transform 1 0 67804 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_728
timestamp 1704896540
transform 1 0 67988 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_740
timestamp 1704896540
transform 1 0 69092 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_752
timestamp 1704896540
transform 1 0 70196 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_764
timestamp 1704896540
transform 1 0 71300 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_776
timestamp 1704896540
transform 1 0 72404 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_782
timestamp 1704896540
transform 1 0 72956 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_784
timestamp 1704896540
transform 1 0 73140 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72_796
timestamp 1704896540
transform 1 0 74244 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_800
timestamp 1704896540
transform 1 0 74612 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_702
timestamp 1704896540
transform 1 0 65596 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_706
timestamp 1704896540
transform 1 0 65964 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_718
timestamp 1704896540
transform 1 0 67068 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_730
timestamp 1704896540
transform 1 0 68172 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_742
timestamp 1704896540
transform 1 0 69276 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_754
timestamp 1704896540
transform 1 0 70380 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_756
timestamp 1704896540
transform 1 0 70564 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_768
timestamp 1704896540
transform 1 0 71668 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_780
timestamp 1704896540
transform 1 0 72772 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73_792
timestamp 1704896540
transform 1 0 73876 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_800
timestamp 1704896540
transform 1 0 74612 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_702
timestamp 1704896540
transform 1 0 65596 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_74_722
timestamp 1704896540
transform 1 0 67436 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_726
timestamp 1704896540
transform 1 0 67804 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_728
timestamp 1704896540
transform 1 0 67988 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_740
timestamp 1704896540
transform 1 0 69092 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_752
timestamp 1704896540
transform 1 0 70196 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_764
timestamp 1704896540
transform 1 0 71300 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_776
timestamp 1704896540
transform 1 0 72404 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_782
timestamp 1704896540
transform 1 0 72956 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_784
timestamp 1704896540
transform 1 0 73140 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_74_796
timestamp 1704896540
transform 1 0 74244 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_800
timestamp 1704896540
transform 1 0 74612 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_710
timestamp 1704896540
transform 1 0 66332 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_722
timestamp 1704896540
transform 1 0 67436 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_734
timestamp 1704896540
transform 1 0 68540 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_75_746
timestamp 1704896540
transform 1 0 69644 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_754
timestamp 1704896540
transform 1 0 70380 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_756
timestamp 1704896540
transform 1 0 70564 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_768
timestamp 1704896540
transform 1 0 71668 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_780
timestamp 1704896540
transform 1 0 72772 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_75_792
timestamp 1704896540
transform 1 0 73876 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_800
timestamp 1704896540
transform 1 0 74612 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_705
timestamp 1704896540
transform 1 0 65872 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_76_717
timestamp 1704896540
transform 1 0 66976 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76_725
timestamp 1704896540
transform 1 0 67712 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_736
timestamp 1704896540
transform 1 0 68724 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_748
timestamp 1704896540
transform 1 0 69828 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_760
timestamp 1704896540
transform 1 0 70932 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_76_772
timestamp 1704896540
transform 1 0 72036 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_76_780
timestamp 1704896540
transform 1 0 72772 0 1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_784
timestamp 1704896540
transform 1 0 73140 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_76_796
timestamp 1704896540
transform 1 0 74244 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_800
timestamp 1704896540
transform 1 0 74612 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_702
timestamp 1704896540
transform 1 0 65596 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_714
timestamp 1704896540
transform 1 0 66700 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_726
timestamp 1704896540
transform 1 0 67804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_738
timestamp 1704896540
transform 1 0 68908 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_77_750
timestamp 1704896540
transform 1 0 70012 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_754
timestamp 1704896540
transform 1 0 70380 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_756
timestamp 1704896540
transform 1 0 70564 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_768
timestamp 1704896540
transform 1 0 71668 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_780
timestamp 1704896540
transform 1 0 72772 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_77_792
timestamp 1704896540
transform 1 0 73876 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_800
timestamp 1704896540
transform 1 0 74612 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_713
timestamp 1704896540
transform 1 0 66608 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_78_725
timestamp 1704896540
transform 1 0 67712 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_728
timestamp 1704896540
transform 1 0 67988 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_740
timestamp 1704896540
transform 1 0 69092 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_752
timestamp 1704896540
transform 1 0 70196 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_764
timestamp 1704896540
transform 1 0 71300 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_776
timestamp 1704896540
transform 1 0 72404 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_782
timestamp 1704896540
transform 1 0 72956 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_784
timestamp 1704896540
transform 1 0 73140 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_78_796
timestamp 1704896540
transform 1 0 74244 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_800
timestamp 1704896540
transform 1 0 74612 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_702
timestamp 1704896540
transform 1 0 65596 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_714
timestamp 1704896540
transform 1 0 66700 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_726
timestamp 1704896540
transform 1 0 67804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_738
timestamp 1704896540
transform 1 0 68908 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_79_750
timestamp 1704896540
transform 1 0 70012 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_754
timestamp 1704896540
transform 1 0 70380 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_756
timestamp 1704896540
transform 1 0 70564 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_768
timestamp 1704896540
transform 1 0 71668 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_780
timestamp 1704896540
transform 1 0 72772 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_79_792
timestamp 1704896540
transform 1 0 73876 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_800
timestamp 1704896540
transform 1 0 74612 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_702
timestamp 1704896540
transform 1 0 65596 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_714
timestamp 1704896540
transform 1 0 66700 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_726
timestamp 1704896540
transform 1 0 67804 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_728
timestamp 1704896540
transform 1 0 67988 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_740
timestamp 1704896540
transform 1 0 69092 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_752
timestamp 1704896540
transform 1 0 70196 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_764
timestamp 1704896540
transform 1 0 71300 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_776
timestamp 1704896540
transform 1 0 72404 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_782
timestamp 1704896540
transform 1 0 72956 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_784
timestamp 1704896540
transform 1 0 73140 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80_796
timestamp 1704896540
transform 1 0 74244 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_800
timestamp 1704896540
transform 1 0 74612 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_710
timestamp 1704896540
transform 1 0 66332 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_722
timestamp 1704896540
transform 1 0 67436 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_734
timestamp 1704896540
transform 1 0 68540 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_81_746
timestamp 1704896540
transform 1 0 69644 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_754
timestamp 1704896540
transform 1 0 70380 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_756
timestamp 1704896540
transform 1 0 70564 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_768
timestamp 1704896540
transform 1 0 71668 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_780
timestamp 1704896540
transform 1 0 72772 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_81_792
timestamp 1704896540
transform 1 0 73876 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_800
timestamp 1704896540
transform 1 0 74612 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_702
timestamp 1704896540
transform 1 0 65596 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_714
timestamp 1704896540
transform 1 0 66700 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_726
timestamp 1704896540
transform 1 0 67804 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_728
timestamp 1704896540
transform 1 0 67988 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_740
timestamp 1704896540
transform 1 0 69092 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_752
timestamp 1704896540
transform 1 0 70196 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_764
timestamp 1704896540
transform 1 0 71300 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_776
timestamp 1704896540
transform 1 0 72404 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_782
timestamp 1704896540
transform 1 0 72956 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_784
timestamp 1704896540
transform 1 0 73140 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_82_796
timestamp 1704896540
transform 1 0 74244 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_800
timestamp 1704896540
transform 1 0 74612 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_702
timestamp 1704896540
transform 1 0 65596 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_714
timestamp 1704896540
transform 1 0 66700 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_726
timestamp 1704896540
transform 1 0 67804 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_738
timestamp 1704896540
transform 1 0 68908 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_83_750
timestamp 1704896540
transform 1 0 70012 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_754
timestamp 1704896540
transform 1 0 70380 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_756
timestamp 1704896540
transform 1 0 70564 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_768
timestamp 1704896540
transform 1 0 71668 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_780
timestamp 1704896540
transform 1 0 72772 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_83_792
timestamp 1704896540
transform 1 0 73876 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_800
timestamp 1704896540
transform 1 0 74612 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_84_716
timestamp 1704896540
transform 1 0 66884 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_84_724
timestamp 1704896540
transform 1 0 67620 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_728
timestamp 1704896540
transform 1 0 67988 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_740
timestamp 1704896540
transform 1 0 69092 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_752
timestamp 1704896540
transform 1 0 70196 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_764
timestamp 1704896540
transform 1 0 71300 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_776
timestamp 1704896540
transform 1 0 72404 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_782
timestamp 1704896540
transform 1 0 72956 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_784
timestamp 1704896540
transform 1 0 73140 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_84_796
timestamp 1704896540
transform 1 0 74244 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_800
timestamp 1704896540
transform 1 0 74612 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_702
timestamp 1704896540
transform 1 0 65596 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_714
timestamp 1704896540
transform 1 0 66700 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_726
timestamp 1704896540
transform 1 0 67804 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_738
timestamp 1704896540
transform 1 0 68908 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85_750
timestamp 1704896540
transform 1 0 70012 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_754
timestamp 1704896540
transform 1 0 70380 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_756
timestamp 1704896540
transform 1 0 70564 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_768
timestamp 1704896540
transform 1 0 71668 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_780
timestamp 1704896540
transform 1 0 72772 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85_792
timestamp 1704896540
transform 1 0 73876 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_800
timestamp 1704896540
transform 1 0 74612 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_702
timestamp 1704896540
transform 1 0 65596 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_714
timestamp 1704896540
transform 1 0 66700 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_726
timestamp 1704896540
transform 1 0 67804 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_728
timestamp 1704896540
transform 1 0 67988 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_740
timestamp 1704896540
transform 1 0 69092 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_752
timestamp 1704896540
transform 1 0 70196 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_764
timestamp 1704896540
transform 1 0 71300 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_776
timestamp 1704896540
transform 1 0 72404 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_782
timestamp 1704896540
transform 1 0 72956 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_784
timestamp 1704896540
transform 1 0 73140 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_86_796
timestamp 1704896540
transform 1 0 74244 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_800
timestamp 1704896540
transform 1 0 74612 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_710
timestamp 1704896540
transform 1 0 66332 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_722
timestamp 1704896540
transform 1 0 67436 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_734
timestamp 1704896540
transform 1 0 68540 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_87_746
timestamp 1704896540
transform 1 0 69644 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_754
timestamp 1704896540
transform 1 0 70380 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_756
timestamp 1704896540
transform 1 0 70564 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_768
timestamp 1704896540
transform 1 0 71668 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_780
timestamp 1704896540
transform 1 0 72772 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_87_792
timestamp 1704896540
transform 1 0 73876 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_800
timestamp 1704896540
transform 1 0 74612 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_705
timestamp 1704896540
transform 1 0 65872 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_88_717
timestamp 1704896540
transform 1 0 66976 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_88_725
timestamp 1704896540
transform 1 0 67712 0 1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_728
timestamp 1704896540
transform 1 0 67988 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_740
timestamp 1704896540
transform 1 0 69092 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_752
timestamp 1704896540
transform 1 0 70196 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_764
timestamp 1704896540
transform 1 0 71300 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_776
timestamp 1704896540
transform 1 0 72404 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_782
timestamp 1704896540
transform 1 0 72956 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_784
timestamp 1704896540
transform 1 0 73140 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_88_796
timestamp 1704896540
transform 1 0 74244 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_800
timestamp 1704896540
transform 1 0 74612 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_705
timestamp 1704896540
transform 1 0 65872 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_717
timestamp 1704896540
transform 1 0 66976 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_729
timestamp 1704896540
transform 1 0 68080 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_741
timestamp 1704896540
transform 1 0 69184 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_89_753
timestamp 1704896540
transform 1 0 70288 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_756
timestamp 1704896540
transform 1 0 70564 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_768
timestamp 1704896540
transform 1 0 71668 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_780
timestamp 1704896540
transform 1 0 72772 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_89_792
timestamp 1704896540
transform 1 0 73876 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_800
timestamp 1704896540
transform 1 0 74612 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_713
timestamp 1704896540
transform 1 0 66608 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_90_725
timestamp 1704896540
transform 1 0 67712 0 1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_728
timestamp 1704896540
transform 1 0 67988 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_740
timestamp 1704896540
transform 1 0 69092 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_752
timestamp 1704896540
transform 1 0 70196 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_764
timestamp 1704896540
transform 1 0 71300 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_776
timestamp 1704896540
transform 1 0 72404 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_782
timestamp 1704896540
transform 1 0 72956 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_784
timestamp 1704896540
transform 1 0 73140 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_90_796
timestamp 1704896540
transform 1 0 74244 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_800
timestamp 1704896540
transform 1 0 74612 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_702
timestamp 1704896540
transform 1 0 65596 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_714
timestamp 1704896540
transform 1 0 66700 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_726
timestamp 1704896540
transform 1 0 67804 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_738
timestamp 1704896540
transform 1 0 68908 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_91_750
timestamp 1704896540
transform 1 0 70012 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_754
timestamp 1704896540
transform 1 0 70380 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_756
timestamp 1704896540
transform 1 0 70564 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_768
timestamp 1704896540
transform 1 0 71668 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_780
timestamp 1704896540
transform 1 0 72772 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_91_792
timestamp 1704896540
transform 1 0 73876 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_800
timestamp 1704896540
transform 1 0 74612 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_702
timestamp 1704896540
transform 1 0 65596 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_714
timestamp 1704896540
transform 1 0 66700 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_726
timestamp 1704896540
transform 1 0 67804 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_728
timestamp 1704896540
transform 1 0 67988 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_740
timestamp 1704896540
transform 1 0 69092 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_752
timestamp 1704896540
transform 1 0 70196 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_764
timestamp 1704896540
transform 1 0 71300 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_776
timestamp 1704896540
transform 1 0 72404 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_782
timestamp 1704896540
transform 1 0 72956 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_784
timestamp 1704896540
transform 1 0 73140 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_92_796
timestamp 1704896540
transform 1 0 74244 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_800
timestamp 1704896540
transform 1 0 74612 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_710
timestamp 1704896540
transform 1 0 66332 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_722
timestamp 1704896540
transform 1 0 67436 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_734
timestamp 1704896540
transform 1 0 68540 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_93_746
timestamp 1704896540
transform 1 0 69644 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_754
timestamp 1704896540
transform 1 0 70380 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_756
timestamp 1704896540
transform 1 0 70564 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_768
timestamp 1704896540
transform 1 0 71668 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_780
timestamp 1704896540
transform 1 0 72772 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_93_792
timestamp 1704896540
transform 1 0 73876 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_800
timestamp 1704896540
transform 1 0 74612 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_708
timestamp 1704896540
transform 1 0 66148 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_720
timestamp 1704896540
transform 1 0 67252 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_726
timestamp 1704896540
transform 1 0 67804 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_728
timestamp 1704896540
transform 1 0 67988 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_740
timestamp 1704896540
transform 1 0 69092 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_752
timestamp 1704896540
transform 1 0 70196 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_764
timestamp 1704896540
transform 1 0 71300 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_776
timestamp 1704896540
transform 1 0 72404 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_782
timestamp 1704896540
transform 1 0 72956 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_784
timestamp 1704896540
transform 1 0 73140 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_94_796
timestamp 1704896540
transform 1 0 74244 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_800
timestamp 1704896540
transform 1 0 74612 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_710
timestamp 1704896540
transform 1 0 66332 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_722
timestamp 1704896540
transform 1 0 67436 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_734
timestamp 1704896540
transform 1 0 68540 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_95_746
timestamp 1704896540
transform 1 0 69644 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_754
timestamp 1704896540
transform 1 0 70380 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_756
timestamp 1704896540
transform 1 0 70564 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_768
timestamp 1704896540
transform 1 0 71668 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_780
timestamp 1704896540
transform 1 0 72772 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_95_792
timestamp 1704896540
transform 1 0 73876 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_800
timestamp 1704896540
transform 1 0 74612 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_96_718
timestamp 1704896540
transform 1 0 67068 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_726
timestamp 1704896540
transform 1 0 67804 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_728
timestamp 1704896540
transform 1 0 67988 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_740
timestamp 1704896540
transform 1 0 69092 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_752
timestamp 1704896540
transform 1 0 70196 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_764
timestamp 1704896540
transform 1 0 71300 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_776
timestamp 1704896540
transform 1 0 72404 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_782
timestamp 1704896540
transform 1 0 72956 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_784
timestamp 1704896540
transform 1 0 73140 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_96_796
timestamp 1704896540
transform 1 0 74244 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_800
timestamp 1704896540
transform 1 0 74612 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_702
timestamp 1704896540
transform 1 0 65596 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_714
timestamp 1704896540
transform 1 0 66700 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_726
timestamp 1704896540
transform 1 0 67804 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_738
timestamp 1704896540
transform 1 0 68908 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_97_750
timestamp 1704896540
transform 1 0 70012 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_754
timestamp 1704896540
transform 1 0 70380 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_756
timestamp 1704896540
transform 1 0 70564 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_768
timestamp 1704896540
transform 1 0 71668 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_780
timestamp 1704896540
transform 1 0 72772 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_97_792
timestamp 1704896540
transform 1 0 73876 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_800
timestamp 1704896540
transform 1 0 74612 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_702
timestamp 1704896540
transform 1 0 65596 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_714
timestamp 1704896540
transform 1 0 66700 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_726
timestamp 1704896540
transform 1 0 67804 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_728
timestamp 1704896540
transform 1 0 67988 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_740
timestamp 1704896540
transform 1 0 69092 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_752
timestamp 1704896540
transform 1 0 70196 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_764
timestamp 1704896540
transform 1 0 71300 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_776
timestamp 1704896540
transform 1 0 72404 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_782
timestamp 1704896540
transform 1 0 72956 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_784
timestamp 1704896540
transform 1 0 73140 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_98_796
timestamp 1704896540
transform 1 0 74244 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_800
timestamp 1704896540
transform 1 0 74612 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_710
timestamp 1704896540
transform 1 0 66332 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_722
timestamp 1704896540
transform 1 0 67436 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_734
timestamp 1704896540
transform 1 0 68540 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_99_746
timestamp 1704896540
transform 1 0 69644 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_754
timestamp 1704896540
transform 1 0 70380 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_756
timestamp 1704896540
transform 1 0 70564 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_768
timestamp 1704896540
transform 1 0 71668 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_780
timestamp 1704896540
transform 1 0 72772 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_99_792
timestamp 1704896540
transform 1 0 73876 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_800
timestamp 1704896540
transform 1 0 74612 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_702
timestamp 1704896540
transform 1 0 65596 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_714
timestamp 1704896540
transform 1 0 66700 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_726
timestamp 1704896540
transform 1 0 67804 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_728
timestamp 1704896540
transform 1 0 67988 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_740
timestamp 1704896540
transform 1 0 69092 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_752
timestamp 1704896540
transform 1 0 70196 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_764
timestamp 1704896540
transform 1 0 71300 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_776
timestamp 1704896540
transform 1 0 72404 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_782
timestamp 1704896540
transform 1 0 72956 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_784
timestamp 1704896540
transform 1 0 73140 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_100_796
timestamp 1704896540
transform 1 0 74244 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_800
timestamp 1704896540
transform 1 0 74612 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_702
timestamp 1704896540
transform 1 0 65596 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_714
timestamp 1704896540
transform 1 0 66700 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_726
timestamp 1704896540
transform 1 0 67804 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_738
timestamp 1704896540
transform 1 0 68908 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_101_750
timestamp 1704896540
transform 1 0 70012 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_754
timestamp 1704896540
transform 1 0 70380 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_756
timestamp 1704896540
transform 1 0 70564 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_768
timestamp 1704896540
transform 1 0 71668 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_780
timestamp 1704896540
transform 1 0 72772 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_101_792
timestamp 1704896540
transform 1 0 73876 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_800
timestamp 1704896540
transform 1 0 74612 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_710
timestamp 1704896540
transform 1 0 66332 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_102_722
timestamp 1704896540
transform 1 0 67436 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_726
timestamp 1704896540
transform 1 0 67804 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_728
timestamp 1704896540
transform 1 0 67988 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_740
timestamp 1704896540
transform 1 0 69092 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_752
timestamp 1704896540
transform 1 0 70196 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_764
timestamp 1704896540
transform 1 0 71300 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_102_776
timestamp 1704896540
transform 1 0 72404 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_782
timestamp 1704896540
transform 1 0 72956 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_784
timestamp 1704896540
transform 1 0 73140 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_102_796
timestamp 1704896540
transform 1 0 74244 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_800
timestamp 1704896540
transform 1 0 74612 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_702
timestamp 1704896540
transform 1 0 65596 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_714
timestamp 1704896540
transform 1 0 66700 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_726
timestamp 1704896540
transform 1 0 67804 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_738
timestamp 1704896540
transform 1 0 68908 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_103_750
timestamp 1704896540
transform 1 0 70012 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103_754
timestamp 1704896540
transform 1 0 70380 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_756
timestamp 1704896540
transform 1 0 70564 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_768
timestamp 1704896540
transform 1 0 71668 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_780
timestamp 1704896540
transform 1 0 72772 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_103_792
timestamp 1704896540
transform 1 0 73876 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103_800
timestamp 1704896540
transform 1 0 74612 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_702
timestamp 1704896540
transform 1 0 65596 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_714
timestamp 1704896540
transform 1 0 66700 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_726
timestamp 1704896540
transform 1 0 67804 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_728
timestamp 1704896540
transform 1 0 67988 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_740
timestamp 1704896540
transform 1 0 69092 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_752
timestamp 1704896540
transform 1 0 70196 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_764
timestamp 1704896540
transform 1 0 71300 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_104_776
timestamp 1704896540
transform 1 0 72404 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_782
timestamp 1704896540
transform 1 0 72956 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_784
timestamp 1704896540
transform 1 0 73140 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_104_796
timestamp 1704896540
transform 1 0 74244 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_800
timestamp 1704896540
transform 1 0 74612 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_710
timestamp 1704896540
transform 1 0 66332 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_722
timestamp 1704896540
transform 1 0 67436 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_734
timestamp 1704896540
transform 1 0 68540 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_105_746
timestamp 1704896540
transform 1 0 69644 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_105_754
timestamp 1704896540
transform 1 0 70380 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_756
timestamp 1704896540
transform 1 0 70564 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_768
timestamp 1704896540
transform 1 0 71668 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_780
timestamp 1704896540
transform 1 0 72772 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_105_792
timestamp 1704896540
transform 1 0 73876 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_105_800
timestamp 1704896540
transform 1 0 74612 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_702
timestamp 1704896540
transform 1 0 65596 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_714
timestamp 1704896540
transform 1 0 66700 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_726
timestamp 1704896540
transform 1 0 67804 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_728
timestamp 1704896540
transform 1 0 67988 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_740
timestamp 1704896540
transform 1 0 69092 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_752
timestamp 1704896540
transform 1 0 70196 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_764
timestamp 1704896540
transform 1 0 71300 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106_776
timestamp 1704896540
transform 1 0 72404 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_782
timestamp 1704896540
transform 1 0 72956 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_784
timestamp 1704896540
transform 1 0 73140 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_106_796
timestamp 1704896540
transform 1 0 74244 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_800
timestamp 1704896540
transform 1 0 74612 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_702
timestamp 1704896540
transform 1 0 65596 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_714
timestamp 1704896540
transform 1 0 66700 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_726
timestamp 1704896540
transform 1 0 67804 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_738
timestamp 1704896540
transform 1 0 68908 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_107_750
timestamp 1704896540
transform 1 0 70012 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_107_754
timestamp 1704896540
transform 1 0 70380 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_756
timestamp 1704896540
transform 1 0 70564 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_768
timestamp 1704896540
transform 1 0 71668 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_780
timestamp 1704896540
transform 1 0 72772 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_107_792
timestamp 1704896540
transform 1 0 73876 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_107_800
timestamp 1704896540
transform 1 0 74612 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_710
timestamp 1704896540
transform 1 0 66332 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_108_722
timestamp 1704896540
transform 1 0 67436 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_726
timestamp 1704896540
transform 1 0 67804 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_728
timestamp 1704896540
transform 1 0 67988 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_740
timestamp 1704896540
transform 1 0 69092 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_752
timestamp 1704896540
transform 1 0 70196 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_764
timestamp 1704896540
transform 1 0 71300 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_108_776
timestamp 1704896540
transform 1 0 72404 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_782
timestamp 1704896540
transform 1 0 72956 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_784
timestamp 1704896540
transform 1 0 73140 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_108_796
timestamp 1704896540
transform 1 0 74244 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_800
timestamp 1704896540
transform 1 0 74612 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_702
timestamp 1704896540
transform 1 0 65596 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_714
timestamp 1704896540
transform 1 0 66700 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_726
timestamp 1704896540
transform 1 0 67804 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_738
timestamp 1704896540
transform 1 0 68908 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_109_750
timestamp 1704896540
transform 1 0 70012 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_109_754
timestamp 1704896540
transform 1 0 70380 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_756
timestamp 1704896540
transform 1 0 70564 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_768
timestamp 1704896540
transform 1 0 71668 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_780
timestamp 1704896540
transform 1 0 72772 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_109_792
timestamp 1704896540
transform 1 0 73876 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_109_800
timestamp 1704896540
transform 1 0 74612 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_702
timestamp 1704896540
transform 1 0 65596 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_714
timestamp 1704896540
transform 1 0 66700 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_726
timestamp 1704896540
transform 1 0 67804 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_728
timestamp 1704896540
transform 1 0 67988 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_740
timestamp 1704896540
transform 1 0 69092 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_752
timestamp 1704896540
transform 1 0 70196 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_764
timestamp 1704896540
transform 1 0 71300 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_110_776
timestamp 1704896540
transform 1 0 72404 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_782
timestamp 1704896540
transform 1 0 72956 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_784
timestamp 1704896540
transform 1 0 73140 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_110_796
timestamp 1704896540
transform 1 0 74244 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_800
timestamp 1704896540
transform 1 0 74612 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_710
timestamp 1704896540
transform 1 0 66332 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_722
timestamp 1704896540
transform 1 0 67436 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_734
timestamp 1704896540
transform 1 0 68540 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_111_746
timestamp 1704896540
transform 1 0 69644 0 -1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111_754
timestamp 1704896540
transform 1 0 70380 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_756
timestamp 1704896540
transform 1 0 70564 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_768
timestamp 1704896540
transform 1 0 71668 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_780
timestamp 1704896540
transform 1 0 72772 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_111_792
timestamp 1704896540
transform 1 0 73876 0 -1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111_800
timestamp 1704896540
transform 1 0 74612 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_702
timestamp 1704896540
transform 1 0 65596 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_714
timestamp 1704896540
transform 1 0 66700 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112_726
timestamp 1704896540
transform 1 0 67804 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_728
timestamp 1704896540
transform 1 0 67988 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_740
timestamp 1704896540
transform 1 0 69092 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_752
timestamp 1704896540
transform 1 0 70196 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_764
timestamp 1704896540
transform 1 0 71300 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_112_776
timestamp 1704896540
transform 1 0 72404 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112_782
timestamp 1704896540
transform 1 0 72956 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_784
timestamp 1704896540
transform 1 0 73140 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_112_796
timestamp 1704896540
transform 1 0 74244 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112_800
timestamp 1704896540
transform 1 0 74612 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_702
timestamp 1704896540
transform 1 0 65596 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_714
timestamp 1704896540
transform 1 0 66700 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_726
timestamp 1704896540
transform 1 0 67804 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_738
timestamp 1704896540
transform 1 0 68908 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_113_750
timestamp 1704896540
transform 1 0 70012 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113_754
timestamp 1704896540
transform 1 0 70380 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_756
timestamp 1704896540
transform 1 0 70564 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_768
timestamp 1704896540
transform 1 0 71668 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_780
timestamp 1704896540
transform 1 0 72772 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_113_792
timestamp 1704896540
transform 1 0 73876 0 -1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113_800
timestamp 1704896540
transform 1 0 74612 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_702
timestamp 1704896540
transform 1 0 65596 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_711
timestamp 1704896540
transform 1 0 66424 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_114_723
timestamp 1704896540
transform 1 0 67528 0 1 63104
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_728
timestamp 1704896540
transform 1 0 67988 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_740
timestamp 1704896540
transform 1 0 69092 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_752
timestamp 1704896540
transform 1 0 70196 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_764
timestamp 1704896540
transform 1 0 71300 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_114_776
timestamp 1704896540
transform 1 0 72404 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_782
timestamp 1704896540
transform 1 0 72956 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_784
timestamp 1704896540
transform 1 0 73140 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_114_796
timestamp 1704896540
transform 1 0 74244 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_800
timestamp 1704896540
transform 1 0 74612 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_702
timestamp 1704896540
transform 1 0 65596 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_714
timestamp 1704896540
transform 1 0 66700 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_726
timestamp 1704896540
transform 1 0 67804 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_738
timestamp 1704896540
transform 1 0 68908 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_115_750
timestamp 1704896540
transform 1 0 70012 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115_754
timestamp 1704896540
transform 1 0 70380 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_756
timestamp 1704896540
transform 1 0 70564 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_768
timestamp 1704896540
transform 1 0 71668 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_780
timestamp 1704896540
transform 1 0 72772 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_115_792
timestamp 1704896540
transform 1 0 73876 0 -1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115_800
timestamp 1704896540
transform 1 0 74612 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_702
timestamp 1704896540
transform 1 0 65596 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_714
timestamp 1704896540
transform 1 0 66700 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_726
timestamp 1704896540
transform 1 0 67804 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_728
timestamp 1704896540
transform 1 0 67988 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_740
timestamp 1704896540
transform 1 0 69092 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_752
timestamp 1704896540
transform 1 0 70196 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_764
timestamp 1704896540
transform 1 0 71300 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_116_776
timestamp 1704896540
transform 1 0 72404 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_782
timestamp 1704896540
transform 1 0 72956 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_784
timestamp 1704896540
transform 1 0 73140 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_116_796
timestamp 1704896540
transform 1 0 74244 0 1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_800
timestamp 1704896540
transform 1 0 74612 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_702
timestamp 1704896540
transform 1 0 65596 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_714
timestamp 1704896540
transform 1 0 66700 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_726
timestamp 1704896540
transform 1 0 67804 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_738
timestamp 1704896540
transform 1 0 68908 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_117_750
timestamp 1704896540
transform 1 0 70012 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117_754
timestamp 1704896540
transform 1 0 70380 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_756
timestamp 1704896540
transform 1 0 70564 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_768
timestamp 1704896540
transform 1 0 71668 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_780
timestamp 1704896540
transform 1 0 72772 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_117_792
timestamp 1704896540
transform 1 0 73876 0 -1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117_800
timestamp 1704896540
transform 1 0 74612 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_702
timestamp 1704896540
transform 1 0 65596 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_714
timestamp 1704896540
transform 1 0 66700 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_726
timestamp 1704896540
transform 1 0 67804 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_728
timestamp 1704896540
transform 1 0 67988 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_740
timestamp 1704896540
transform 1 0 69092 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_752
timestamp 1704896540
transform 1 0 70196 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_764
timestamp 1704896540
transform 1 0 71300 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118_776
timestamp 1704896540
transform 1 0 72404 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_782
timestamp 1704896540
transform 1 0 72956 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_784
timestamp 1704896540
transform 1 0 73140 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_118_796
timestamp 1704896540
transform 1 0 74244 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_800
timestamp 1704896540
transform 1 0 74612 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_702
timestamp 1704896540
transform 1 0 65596 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_714
timestamp 1704896540
transform 1 0 66700 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_726
timestamp 1704896540
transform 1 0 67804 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_738
timestamp 1704896540
transform 1 0 68908 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_119_750
timestamp 1704896540
transform 1 0 70012 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119_754
timestamp 1704896540
transform 1 0 70380 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_756
timestamp 1704896540
transform 1 0 70564 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_768
timestamp 1704896540
transform 1 0 71668 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_780
timestamp 1704896540
transform 1 0 72772 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_119_792
timestamp 1704896540
transform 1 0 73876 0 -1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119_800
timestamp 1704896540
transform 1 0 74612 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_702
timestamp 1704896540
transform 1 0 65596 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_714
timestamp 1704896540
transform 1 0 66700 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_120_726
timestamp 1704896540
transform 1 0 67804 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_728
timestamp 1704896540
transform 1 0 67988 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_740
timestamp 1704896540
transform 1 0 69092 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_752
timestamp 1704896540
transform 1 0 70196 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_764
timestamp 1704896540
transform 1 0 71300 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_120_776
timestamp 1704896540
transform 1 0 72404 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_120_782
timestamp 1704896540
transform 1 0 72956 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_784
timestamp 1704896540
transform 1 0 73140 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_120_796
timestamp 1704896540
transform 1 0 74244 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_120_800
timestamp 1704896540
transform 1 0 74612 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_702
timestamp 1704896540
transform 1 0 65596 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_714
timestamp 1704896540
transform 1 0 66700 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_726
timestamp 1704896540
transform 1 0 67804 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_738
timestamp 1704896540
transform 1 0 68908 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_121_750
timestamp 1704896540
transform 1 0 70012 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_121_754
timestamp 1704896540
transform 1 0 70380 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_756
timestamp 1704896540
transform 1 0 70564 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_768
timestamp 1704896540
transform 1 0 71668 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_780
timestamp 1704896540
transform 1 0 72772 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_121_792
timestamp 1704896540
transform 1 0 73876 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_121_800
timestamp 1704896540
transform 1 0 74612 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_702
timestamp 1704896540
transform 1 0 65596 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_714
timestamp 1704896540
transform 1 0 66700 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_122_726
timestamp 1704896540
transform 1 0 67804 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_728
timestamp 1704896540
transform 1 0 67988 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_740
timestamp 1704896540
transform 1 0 69092 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_752
timestamp 1704896540
transform 1 0 70196 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_764
timestamp 1704896540
transform 1 0 71300 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_122_776
timestamp 1704896540
transform 1 0 72404 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_122_782
timestamp 1704896540
transform 1 0 72956 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_784
timestamp 1704896540
transform 1 0 73140 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_122_796
timestamp 1704896540
transform 1 0 74244 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_122_800
timestamp 1704896540
transform 1 0 74612 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_702
timestamp 1704896540
transform 1 0 65596 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_714
timestamp 1704896540
transform 1 0 66700 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_726
timestamp 1704896540
transform 1 0 67804 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_738
timestamp 1704896540
transform 1 0 68908 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_123_750
timestamp 1704896540
transform 1 0 70012 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_123_754
timestamp 1704896540
transform 1 0 70380 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_756
timestamp 1704896540
transform 1 0 70564 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_768
timestamp 1704896540
transform 1 0 71668 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_780
timestamp 1704896540
transform 1 0 72772 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_123_792
timestamp 1704896540
transform 1 0 73876 0 -1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_123_800
timestamp 1704896540
transform 1 0 74612 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_124_702
timestamp 1704896540
transform 1 0 65596 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_124_714
timestamp 1704896540
transform 1 0 66700 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_124_726
timestamp 1704896540
transform 1 0 67804 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_124_728
timestamp 1704896540
transform 1 0 67988 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_124_740
timestamp 1704896540
transform 1 0 69092 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_124_752
timestamp 1704896540
transform 1 0 70196 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_124_764
timestamp 1704896540
transform 1 0 71300 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_124_776
timestamp 1704896540
transform 1 0 72404 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_124_782
timestamp 1704896540
transform 1 0 72956 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_124_784
timestamp 1704896540
transform 1 0 73140 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_124_796
timestamp 1704896540
transform 1 0 74244 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_124_800
timestamp 1704896540
transform 1 0 74612 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125_702
timestamp 1704896540
transform 1 0 65596 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125_714
timestamp 1704896540
transform 1 0 66700 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125_726
timestamp 1704896540
transform 1 0 67804 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125_738
timestamp 1704896540
transform 1 0 68908 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_125_750
timestamp 1704896540
transform 1 0 70012 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_125_754
timestamp 1704896540
transform 1 0 70380 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125_756
timestamp 1704896540
transform 1 0 70564 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125_768
timestamp 1704896540
transform 1 0 71668 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125_780
timestamp 1704896540
transform 1 0 72772 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_125_792
timestamp 1704896540
transform 1 0 73876 0 -1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_125_800
timestamp 1704896540
transform 1 0 74612 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_126_702
timestamp 1704896540
transform 1 0 65596 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_126_714
timestamp 1704896540
transform 1 0 66700 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_126_726
timestamp 1704896540
transform 1 0 67804 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_126_728
timestamp 1704896540
transform 1 0 67988 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_126_740
timestamp 1704896540
transform 1 0 69092 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_126_752
timestamp 1704896540
transform 1 0 70196 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_126_764
timestamp 1704896540
transform 1 0 71300 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_126_776
timestamp 1704896540
transform 1 0 72404 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_126_782
timestamp 1704896540
transform 1 0 72956 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_126_784
timestamp 1704896540
transform 1 0 73140 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_126_796
timestamp 1704896540
transform 1 0 74244 0 1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_126_800
timestamp 1704896540
transform 1 0 74612 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_127_702
timestamp 1704896540
transform 1 0 65596 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_127_714
timestamp 1704896540
transform 1 0 66700 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_127_726
timestamp 1704896540
transform 1 0 67804 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_127_738
timestamp 1704896540
transform 1 0 68908 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_127_750
timestamp 1704896540
transform 1 0 70012 0 -1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_127_754
timestamp 1704896540
transform 1 0 70380 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_127_756
timestamp 1704896540
transform 1 0 70564 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_127_768
timestamp 1704896540
transform 1 0 71668 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_127_780
timestamp 1704896540
transform 1 0 72772 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_127_792
timestamp 1704896540
transform 1 0 73876 0 -1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_127_800
timestamp 1704896540
transform 1 0 74612 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_128_702
timestamp 1704896540
transform 1 0 65596 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_128_714
timestamp 1704896540
transform 1 0 66700 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_128_726
timestamp 1704896540
transform 1 0 67804 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_128_728
timestamp 1704896540
transform 1 0 67988 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_128_740
timestamp 1704896540
transform 1 0 69092 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_128_752
timestamp 1704896540
transform 1 0 70196 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_128_764
timestamp 1704896540
transform 1 0 71300 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_128_776
timestamp 1704896540
transform 1 0 72404 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_128_782
timestamp 1704896540
transform 1 0 72956 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_128_784
timestamp 1704896540
transform 1 0 73140 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_128_796
timestamp 1704896540
transform 1 0 74244 0 1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_128_800
timestamp 1704896540
transform 1 0 74612 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_129_702
timestamp 1704896540
transform 1 0 65596 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_129_714
timestamp 1704896540
transform 1 0 66700 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_129_726
timestamp 1704896540
transform 1 0 67804 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_129_738
timestamp 1704896540
transform 1 0 68908 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_129_750
timestamp 1704896540
transform 1 0 70012 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_129_754
timestamp 1704896540
transform 1 0 70380 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_129_756
timestamp 1704896540
transform 1 0 70564 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_129_768
timestamp 1704896540
transform 1 0 71668 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_129_780
timestamp 1704896540
transform 1 0 72772 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_129_792
timestamp 1704896540
transform 1 0 73876 0 -1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_129_800
timestamp 1704896540
transform 1 0 74612 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_130_702
timestamp 1704896540
transform 1 0 65596 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_130_714
timestamp 1704896540
transform 1 0 66700 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_130_726
timestamp 1704896540
transform 1 0 67804 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_130_728
timestamp 1704896540
transform 1 0 67988 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_130_740
timestamp 1704896540
transform 1 0 69092 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_130_752
timestamp 1704896540
transform 1 0 70196 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_130_764
timestamp 1704896540
transform 1 0 71300 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_130_776
timestamp 1704896540
transform 1 0 72404 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_130_782
timestamp 1704896540
transform 1 0 72956 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_130_784
timestamp 1704896540
transform 1 0 73140 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_130_796
timestamp 1704896540
transform 1 0 74244 0 1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_130_800
timestamp 1704896540
transform 1 0 74612 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_131_702
timestamp 1704896540
transform 1 0 65596 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_131_714
timestamp 1704896540
transform 1 0 66700 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_131_726
timestamp 1704896540
transform 1 0 67804 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_131_738
timestamp 1704896540
transform 1 0 68908 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_131_750
timestamp 1704896540
transform 1 0 70012 0 -1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_131_754
timestamp 1704896540
transform 1 0 70380 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_131_756
timestamp 1704896540
transform 1 0 70564 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_131_768
timestamp 1704896540
transform 1 0 71668 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_131_780
timestamp 1704896540
transform 1 0 72772 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_131_792
timestamp 1704896540
transform 1 0 73876 0 -1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_131_800
timestamp 1704896540
transform 1 0 74612 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_132_702
timestamp 1704896540
transform 1 0 65596 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_132_714
timestamp 1704896540
transform 1 0 66700 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_132_726
timestamp 1704896540
transform 1 0 67804 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_132_728
timestamp 1704896540
transform 1 0 67988 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_132_740
timestamp 1704896540
transform 1 0 69092 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_132_752
timestamp 1704896540
transform 1 0 70196 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_132_764
timestamp 1704896540
transform 1 0 71300 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_132_776
timestamp 1704896540
transform 1 0 72404 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_132_782
timestamp 1704896540
transform 1 0 72956 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_132_784
timestamp 1704896540
transform 1 0 73140 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_132_796
timestamp 1704896540
transform 1 0 74244 0 1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_132_800
timestamp 1704896540
transform 1 0 74612 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_133_702
timestamp 1704896540
transform 1 0 65596 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_133_714
timestamp 1704896540
transform 1 0 66700 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_133_726
timestamp 1704896540
transform 1 0 67804 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_133_738
timestamp 1704896540
transform 1 0 68908 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_133_750
timestamp 1704896540
transform 1 0 70012 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_133_754
timestamp 1704896540
transform 1 0 70380 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_133_756
timestamp 1704896540
transform 1 0 70564 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_133_768
timestamp 1704896540
transform 1 0 71668 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_133_780
timestamp 1704896540
transform 1 0 72772 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_133_792
timestamp 1704896540
transform 1 0 73876 0 -1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_133_800
timestamp 1704896540
transform 1 0 74612 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_134_702
timestamp 1704896540
transform 1 0 65596 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_134_714
timestamp 1704896540
transform 1 0 66700 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_134_726
timestamp 1704896540
transform 1 0 67804 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_134_728
timestamp 1704896540
transform 1 0 67988 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_134_740
timestamp 1704896540
transform 1 0 69092 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_134_752
timestamp 1704896540
transform 1 0 70196 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_134_764
timestamp 1704896540
transform 1 0 71300 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_134_776
timestamp 1704896540
transform 1 0 72404 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_134_782
timestamp 1704896540
transform 1 0 72956 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_134_784
timestamp 1704896540
transform 1 0 73140 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_134_796
timestamp 1704896540
transform 1 0 74244 0 1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_134_800
timestamp 1704896540
transform 1 0 74612 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_135_702
timestamp 1704896540
transform 1 0 65596 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_135_714
timestamp 1704896540
transform 1 0 66700 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_135_726
timestamp 1704896540
transform 1 0 67804 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_135_738
timestamp 1704896540
transform 1 0 68908 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_135_750
timestamp 1704896540
transform 1 0 70012 0 -1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_135_754
timestamp 1704896540
transform 1 0 70380 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_135_756
timestamp 1704896540
transform 1 0 70564 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_135_768
timestamp 1704896540
transform 1 0 71668 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_135_780
timestamp 1704896540
transform 1 0 72772 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_135_792
timestamp 1704896540
transform 1 0 73876 0 -1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_135_800
timestamp 1704896540
transform 1 0 74612 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_136_702
timestamp 1704896540
transform 1 0 65596 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_136_714
timestamp 1704896540
transform 1 0 66700 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_136_726
timestamp 1704896540
transform 1 0 67804 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_136_728
timestamp 1704896540
transform 1 0 67988 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_136_740
timestamp 1704896540
transform 1 0 69092 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_136_752
timestamp 1704896540
transform 1 0 70196 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_136_764
timestamp 1704896540
transform 1 0 71300 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_136_776
timestamp 1704896540
transform 1 0 72404 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_136_782
timestamp 1704896540
transform 1 0 72956 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_136_784
timestamp 1704896540
transform 1 0 73140 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_136_796
timestamp 1704896540
transform 1 0 74244 0 1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_136_800
timestamp 1704896540
transform 1 0 74612 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_137_702
timestamp 1704896540
transform 1 0 65596 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_137_714
timestamp 1704896540
transform 1 0 66700 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_137_726
timestamp 1704896540
transform 1 0 67804 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_137_738
timestamp 1704896540
transform 1 0 68908 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_137_750
timestamp 1704896540
transform 1 0 70012 0 -1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_137_754
timestamp 1704896540
transform 1 0 70380 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_137_756
timestamp 1704896540
transform 1 0 70564 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_137_768
timestamp 1704896540
transform 1 0 71668 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_137_780
timestamp 1704896540
transform 1 0 72772 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_137_792
timestamp 1704896540
transform 1 0 73876 0 -1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_137_800
timestamp 1704896540
transform 1 0 74612 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_138_702
timestamp 1704896540
transform 1 0 65596 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_138_714
timestamp 1704896540
transform 1 0 66700 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_138_726
timestamp 1704896540
transform 1 0 67804 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_138_728
timestamp 1704896540
transform 1 0 67988 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_138_740
timestamp 1704896540
transform 1 0 69092 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_138_752
timestamp 1704896540
transform 1 0 70196 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_138_764
timestamp 1704896540
transform 1 0 71300 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_138_776
timestamp 1704896540
transform 1 0 72404 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_138_782
timestamp 1704896540
transform 1 0 72956 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_138_784
timestamp 1704896540
transform 1 0 73140 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_138_796
timestamp 1704896540
transform 1 0 74244 0 1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_138_800
timestamp 1704896540
transform 1 0 74612 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_139_702
timestamp 1704896540
transform 1 0 65596 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_139_714
timestamp 1704896540
transform 1 0 66700 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_139_726
timestamp 1704896540
transform 1 0 67804 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_139_738
timestamp 1704896540
transform 1 0 68908 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_139_750
timestamp 1704896540
transform 1 0 70012 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139_754
timestamp 1704896540
transform 1 0 70380 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_139_756
timestamp 1704896540
transform 1 0 70564 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_139_768
timestamp 1704896540
transform 1 0 71668 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_139_780
timestamp 1704896540
transform 1 0 72772 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_139_792
timestamp 1704896540
transform 1 0 73876 0 -1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139_800
timestamp 1704896540
transform 1 0 74612 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_140_702
timestamp 1704896540
transform 1 0 65596 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_140_714
timestamp 1704896540
transform 1 0 66700 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_140_726
timestamp 1704896540
transform 1 0 67804 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_140_728
timestamp 1704896540
transform 1 0 67988 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_140_740
timestamp 1704896540
transform 1 0 69092 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_140_752
timestamp 1704896540
transform 1 0 70196 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_140_764
timestamp 1704896540
transform 1 0 71300 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_140_776
timestamp 1704896540
transform 1 0 72404 0 1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_140_782
timestamp 1704896540
transform 1 0 72956 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_140_784
timestamp 1704896540
transform 1 0 73140 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_140_796
timestamp 1704896540
transform 1 0 74244 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_140_800
timestamp 1704896540
transform 1 0 74612 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141_702
timestamp 1704896540
transform 1 0 65596 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141_714
timestamp 1704896540
transform 1 0 66700 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141_726
timestamp 1704896540
transform 1 0 67804 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141_738
timestamp 1704896540
transform 1 0 68908 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141_750
timestamp 1704896540
transform 1 0 70012 0 -1 78336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_141_754
timestamp 1704896540
transform 1 0 70380 0 -1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141_756
timestamp 1704896540
transform 1 0 70564 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141_768
timestamp 1704896540
transform 1 0 71668 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141_780
timestamp 1704896540
transform 1 0 72772 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_141_792
timestamp 1704896540
transform 1 0 73876 0 -1 78336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_141_800
timestamp 1704896540
transform 1 0 74612 0 -1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_142_702
timestamp 1704896540
transform 1 0 65596 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_142_714
timestamp 1704896540
transform 1 0 66700 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_142_726
timestamp 1704896540
transform 1 0 67804 0 1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_142_728
timestamp 1704896540
transform 1 0 67988 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_142_740
timestamp 1704896540
transform 1 0 69092 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_142_752
timestamp 1704896540
transform 1 0 70196 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_142_764
timestamp 1704896540
transform 1 0 71300 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_142_776
timestamp 1704896540
transform 1 0 72404 0 1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_142_782
timestamp 1704896540
transform 1 0 72956 0 1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_142_784
timestamp 1704896540
transform 1 0 73140 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_142_796
timestamp 1704896540
transform 1 0 74244 0 1 78336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_142_800
timestamp 1704896540
transform 1 0 74612 0 1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_143_702
timestamp 1704896540
transform 1 0 65596 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_143_714
timestamp 1704896540
transform 1 0 66700 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_143_726
timestamp 1704896540
transform 1 0 67804 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_143_738
timestamp 1704896540
transform 1 0 68908 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_143_750
timestamp 1704896540
transform 1 0 70012 0 -1 79424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_143_754
timestamp 1704896540
transform 1 0 70380 0 -1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_143_756
timestamp 1704896540
transform 1 0 70564 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_143_768
timestamp 1704896540
transform 1 0 71668 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_143_780
timestamp 1704896540
transform 1 0 72772 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_143_792
timestamp 1704896540
transform 1 0 73876 0 -1 79424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_143_800
timestamp 1704896540
transform 1 0 74612 0 -1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_144_702
timestamp 1704896540
transform 1 0 65596 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_144_714
timestamp 1704896540
transform 1 0 66700 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_144_726
timestamp 1704896540
transform 1 0 67804 0 1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_144_728
timestamp 1704896540
transform 1 0 67988 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_144_740
timestamp 1704896540
transform 1 0 69092 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_144_752
timestamp 1704896540
transform 1 0 70196 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_144_764
timestamp 1704896540
transform 1 0 71300 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_144_776
timestamp 1704896540
transform 1 0 72404 0 1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_144_782
timestamp 1704896540
transform 1 0 72956 0 1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_144_784
timestamp 1704896540
transform 1 0 73140 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_144_796
timestamp 1704896540
transform 1 0 74244 0 1 79424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_144_800
timestamp 1704896540
transform 1 0 74612 0 1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_145_702
timestamp 1704896540
transform 1 0 65596 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_145_714
timestamp 1704896540
transform 1 0 66700 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_145_726
timestamp 1704896540
transform 1 0 67804 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_145_738
timestamp 1704896540
transform 1 0 68908 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_145_750
timestamp 1704896540
transform 1 0 70012 0 -1 80512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_145_754
timestamp 1704896540
transform 1 0 70380 0 -1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_145_756
timestamp 1704896540
transform 1 0 70564 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_145_768
timestamp 1704896540
transform 1 0 71668 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_145_780
timestamp 1704896540
transform 1 0 72772 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_145_792
timestamp 1704896540
transform 1 0 73876 0 -1 80512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_145_800
timestamp 1704896540
transform 1 0 74612 0 -1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_146_702
timestamp 1704896540
transform 1 0 65596 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_146_714
timestamp 1704896540
transform 1 0 66700 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_146_726
timestamp 1704896540
transform 1 0 67804 0 1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_146_728
timestamp 1704896540
transform 1 0 67988 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_146_740
timestamp 1704896540
transform 1 0 69092 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_146_752
timestamp 1704896540
transform 1 0 70196 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_146_764
timestamp 1704896540
transform 1 0 71300 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_146_776
timestamp 1704896540
transform 1 0 72404 0 1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_146_782
timestamp 1704896540
transform 1 0 72956 0 1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_146_784
timestamp 1704896540
transform 1 0 73140 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_146_796
timestamp 1704896540
transform 1 0 74244 0 1 80512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_146_800
timestamp 1704896540
transform 1 0 74612 0 1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_147_702
timestamp 1704896540
transform 1 0 65596 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_147_714
timestamp 1704896540
transform 1 0 66700 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_147_726
timestamp 1704896540
transform 1 0 67804 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_147_738
timestamp 1704896540
transform 1 0 68908 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_147_750
timestamp 1704896540
transform 1 0 70012 0 -1 81600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_147_754
timestamp 1704896540
transform 1 0 70380 0 -1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_147_756
timestamp 1704896540
transform 1 0 70564 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_147_768
timestamp 1704896540
transform 1 0 71668 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_147_780
timestamp 1704896540
transform 1 0 72772 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_147_792
timestamp 1704896540
transform 1 0 73876 0 -1 81600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_147_800
timestamp 1704896540
transform 1 0 74612 0 -1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_148_702
timestamp 1704896540
transform 1 0 65596 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_148_714
timestamp 1704896540
transform 1 0 66700 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_148_726
timestamp 1704896540
transform 1 0 67804 0 1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_148_728
timestamp 1704896540
transform 1 0 67988 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_148_740
timestamp 1704896540
transform 1 0 69092 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_148_752
timestamp 1704896540
transform 1 0 70196 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_148_764
timestamp 1704896540
transform 1 0 71300 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_148_776
timestamp 1704896540
transform 1 0 72404 0 1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_148_782
timestamp 1704896540
transform 1 0 72956 0 1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_148_784
timestamp 1704896540
transform 1 0 73140 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_148_796
timestamp 1704896540
transform 1 0 74244 0 1 81600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_148_800
timestamp 1704896540
transform 1 0 74612 0 1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_149_702
timestamp 1704896540
transform 1 0 65596 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_149_714
timestamp 1704896540
transform 1 0 66700 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_149_726
timestamp 1704896540
transform 1 0 67804 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_149_738
timestamp 1704896540
transform 1 0 68908 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_149_750
timestamp 1704896540
transform 1 0 70012 0 -1 82688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_149_754
timestamp 1704896540
transform 1 0 70380 0 -1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_149_756
timestamp 1704896540
transform 1 0 70564 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_149_768
timestamp 1704896540
transform 1 0 71668 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_149_780
timestamp 1704896540
transform 1 0 72772 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_149_792
timestamp 1704896540
transform 1 0 73876 0 -1 82688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_149_800
timestamp 1704896540
transform 1 0 74612 0 -1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_150_702
timestamp 1704896540
transform 1 0 65596 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_150_714
timestamp 1704896540
transform 1 0 66700 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_150_726
timestamp 1704896540
transform 1 0 67804 0 1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_150_728
timestamp 1704896540
transform 1 0 67988 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_150_740
timestamp 1704896540
transform 1 0 69092 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_150_752
timestamp 1704896540
transform 1 0 70196 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_150_764
timestamp 1704896540
transform 1 0 71300 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_150_776
timestamp 1704896540
transform 1 0 72404 0 1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_150_782
timestamp 1704896540
transform 1 0 72956 0 1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_150_784
timestamp 1704896540
transform 1 0 73140 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_150_796
timestamp 1704896540
transform 1 0 74244 0 1 82688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_150_800
timestamp 1704896540
transform 1 0 74612 0 1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_151_702
timestamp 1704896540
transform 1 0 65596 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_151_714
timestamp 1704896540
transform 1 0 66700 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_151_726
timestamp 1704896540
transform 1 0 67804 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_151_738
timestamp 1704896540
transform 1 0 68908 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_151_750
timestamp 1704896540
transform 1 0 70012 0 -1 83776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_151_754
timestamp 1704896540
transform 1 0 70380 0 -1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_151_756
timestamp 1704896540
transform 1 0 70564 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_151_768
timestamp 1704896540
transform 1 0 71668 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_151_780
timestamp 1704896540
transform 1 0 72772 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_151_792
timestamp 1704896540
transform 1 0 73876 0 -1 83776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_151_800
timestamp 1704896540
transform 1 0 74612 0 -1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_152_702
timestamp 1704896540
transform 1 0 65596 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_152_714
timestamp 1704896540
transform 1 0 66700 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_152_726
timestamp 1704896540
transform 1 0 67804 0 1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_152_728
timestamp 1704896540
transform 1 0 67988 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_152_740
timestamp 1704896540
transform 1 0 69092 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_152_752
timestamp 1704896540
transform 1 0 70196 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_152_764
timestamp 1704896540
transform 1 0 71300 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_152_776
timestamp 1704896540
transform 1 0 72404 0 1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_152_782
timestamp 1704896540
transform 1 0 72956 0 1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_152_784
timestamp 1704896540
transform 1 0 73140 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_152_796
timestamp 1704896540
transform 1 0 74244 0 1 83776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_152_800
timestamp 1704896540
transform 1 0 74612 0 1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153_702
timestamp 1704896540
transform 1 0 65596 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153_714
timestamp 1704896540
transform 1 0 66700 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153_726
timestamp 1704896540
transform 1 0 67804 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153_738
timestamp 1704896540
transform 1 0 68908 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_153_750
timestamp 1704896540
transform 1 0 70012 0 -1 84864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_153_754
timestamp 1704896540
transform 1 0 70380 0 -1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153_756
timestamp 1704896540
transform 1 0 70564 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153_768
timestamp 1704896540
transform 1 0 71668 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153_780
timestamp 1704896540
transform 1 0 72772 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_153_792
timestamp 1704896540
transform 1 0 73876 0 -1 84864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_153_800
timestamp 1704896540
transform 1 0 74612 0 -1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_154_702
timestamp 1704896540
transform 1 0 65596 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_154_714
timestamp 1704896540
transform 1 0 66700 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_154_726
timestamp 1704896540
transform 1 0 67804 0 1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_154_728
timestamp 1704896540
transform 1 0 67988 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_154_740
timestamp 1704896540
transform 1 0 69092 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_154_752
timestamp 1704896540
transform 1 0 70196 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_154_764
timestamp 1704896540
transform 1 0 71300 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_154_776
timestamp 1704896540
transform 1 0 72404 0 1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_154_782
timestamp 1704896540
transform 1 0 72956 0 1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_154_784
timestamp 1704896540
transform 1 0 73140 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_154_796
timestamp 1704896540
transform 1 0 74244 0 1 84864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_154_800
timestamp 1704896540
transform 1 0 74612 0 1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_155_702
timestamp 1704896540
transform 1 0 65596 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_155_714
timestamp 1704896540
transform 1 0 66700 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_155_726
timestamp 1704896540
transform 1 0 67804 0 -1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_155_728
timestamp 1704896540
transform 1 0 67988 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_155_740
timestamp 1704896540
transform 1 0 69092 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_155_752
timestamp 1704896540
transform 1 0 70196 0 -1 85952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_155_756
timestamp 1704896540
transform 1 0 70564 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_155_768
timestamp 1704896540
transform 1 0 71668 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_155_780
timestamp 1704896540
transform 1 0 72772 0 -1 85952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_155_784
timestamp 1704896540
transform 1 0 73140 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_155_796
timestamp 1704896540
transform 1 0 74244 0 -1 85952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_155_800
timestamp 1704896540
transform 1 0 74612 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 50416 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1704896540
transform 1 0 56304 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1704896540
transform 1 0 29992 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1704896540
transform 1 0 46644 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1704896540
transform -1 0 46092 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1704896540
transform 1 0 53360 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1704896540
transform -1 0 65320 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1704896540
transform 1 0 65596 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1704896540
transform -1 0 23552 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1704896540
transform 1 0 45448 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1704896540
transform 1 0 42688 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1704896540
transform 1 0 52624 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1704896540
transform 1 0 47840 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1704896540
transform 1 0 56672 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1704896540
transform 1 0 66332 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1704896540
transform -1 0 66332 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1704896540
transform 1 0 20884 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1704896540
transform 1 0 44712 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1704896540
transform -1 0 49312 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1704896540
transform 1 0 55568 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1704896540
transform 1 0 67068 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1704896540
transform -1 0 66332 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1704896540
transform -1 0 40480 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1704896540
transform 1 0 51520 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1704896540
transform 1 0 68908 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1704896540
transform -1 0 67804 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1704896540
transform -1 0 49680 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1704896540
transform 1 0 54832 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1704896540
transform -1 0 72128 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1704896540
transform -1 0 67436 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1704896540
transform 1 0 37260 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1704896540
transform 1 0 50784 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1704896540
transform 1 0 35512 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1704896540
transform 1 0 50048 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1704896540
transform -1 0 47104 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1704896540
transform 1 0 54096 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1704896540
transform 1 0 72128 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 1704896540
transform -1 0 68724 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1704896540
transform 1 0 33028 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 1704896540
transform 1 0 49128 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1704896540
transform 1 0 33028 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1704896540
transform 1 0 48944 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1704896540
transform 1 0 55200 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1704896540
transform 1 0 65596 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 1704896540
transform -1 0 53728 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 1704896540
transform -1 0 67068 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1704896540
transform -1 0 53360 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 1704896540
transform -1 0 66332 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 1704896540
transform 1 0 24564 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold50 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 47472 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 1704896540
transform 1 0 55568 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 1704896540
transform 1 0 65596 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 1704896540
transform 1 0 23552 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 1704896540
transform 1 0 28152 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 1704896540
transform 1 0 38272 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold56
timestamp 1704896540
transform 1 0 55200 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 1704896540
transform 1 0 57408 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp 1704896540
transform 1 0 65596 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 1704896540
transform 1 0 57500 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold60
timestamp 1704896540
transform 1 0 65596 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 1704896540
transform -1 0 24196 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold62
timestamp 1704896540
transform -1 0 27876 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold63
timestamp 1704896540
transform 1 0 26036 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold64
timestamp 1704896540
transform -1 0 31924 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold65
timestamp 1704896540
transform 1 0 47564 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold66
timestamp 1704896540
transform 1 0 61180 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold67
timestamp 1704896540
transform -1 0 66332 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold68
timestamp 1704896540
transform -1 0 62652 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold69
timestamp 1704896540
transform -1 0 67804 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold70
timestamp 1704896540
transform 1 0 62560 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold71
timestamp 1704896540
transform -1 0 68724 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold72
timestamp 1704896540
transform 1 0 63848 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold73
timestamp 1704896540
transform -1 0 67068 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold74
timestamp 1704896540
transform 1 0 21988 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold75
timestamp 1704896540
transform 1 0 45540 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold76
timestamp 1704896540
transform 1 0 23828 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold77
timestamp 1704896540
transform 1 0 25668 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold78
timestamp 1704896540
transform 1 0 37168 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold79
timestamp 1704896540
transform 1 0 65596 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold80
timestamp 1704896540
transform 1 0 22724 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold81
timestamp 1704896540
transform -1 0 26772 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold82
timestamp 1704896540
transform -1 0 28612 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold83
timestamp 1704896540
transform 1 0 27048 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold84
timestamp 1704896540
transform 1 0 65596 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold85
timestamp 1704896540
transform -1 0 31556 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold86
timestamp 1704896540
transform 1 0 31004 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold87
timestamp 1704896540
transform 1 0 39744 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold88
timestamp 1704896540
transform -1 0 67068 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold89
timestamp 1704896540
transform 1 0 26036 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold90
timestamp 1704896540
transform -1 0 27876 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold91
timestamp 1704896540
transform -1 0 32016 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold92
timestamp 1704896540
transform -1 0 33120 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold93
timestamp 1704896540
transform 1 0 65596 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold94
timestamp 1704896540
transform -1 0 33580 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold95
timestamp 1704896540
transform 1 0 32292 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold96
timestamp 1704896540
transform 1 0 41032 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold97
timestamp 1704896540
transform -1 0 67068 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold98
timestamp 1704896540
transform 1 0 30820 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold99
timestamp 1704896540
transform 1 0 30820 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold100
timestamp 1704896540
transform 1 0 31556 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold101
timestamp 1704896540
transform 1 0 44528 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold102
timestamp 1704896540
transform -1 0 67068 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold103
timestamp 1704896540
transform 1 0 41952 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold104
timestamp 1704896540
transform -1 0 66332 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold105
timestamp 1704896540
transform 1 0 40112 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold106
timestamp 1704896540
transform -1 0 67804 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold107
timestamp 1704896540
transform 1 0 38732 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold108
timestamp 1704896540
transform -1 0 67068 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold109
timestamp 1704896540
transform 1 0 35604 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold110
timestamp 1704896540
transform 1 0 66332 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold111
timestamp 1704896540
transform -1 0 34500 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold112
timestamp 1704896540
transform -1 0 66332 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold113
timestamp 1704896540
transform 1 0 35972 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold114
timestamp 1704896540
transform -1 0 66332 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold115
timestamp 1704896540
transform 1 0 30452 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold116
timestamp 1704896540
transform -1 0 66332 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold117
timestamp 1704896540
transform 1 0 28612 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold118
timestamp 1704896540
transform -1 0 66332 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold119
timestamp 1704896540
transform 1 0 29808 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold120
timestamp 1704896540
transform -1 0 66332 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold121
timestamp 1704896540
transform 1 0 23092 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold122
timestamp 1704896540
transform 1 0 29716 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold123
timestamp 1704896540
transform -1 0 66332 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold124
timestamp 1704896540
transform 1 0 20148 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold125
timestamp 1704896540
transform 1 0 25300 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold126
timestamp 1704896540
transform 1 0 33120 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold127
timestamp 1704896540
transform -1 0 66332 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold128
timestamp 1704896540
transform 1 0 22356 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold129
timestamp 1704896540
transform 1 0 26220 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold130
timestamp 1704896540
transform 1 0 27416 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold131
timestamp 1704896540
transform 1 0 27876 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold132
timestamp 1704896540
transform -1 0 25668 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold133
timestamp 1704896540
transform -1 0 25852 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold134
timestamp 1704896540
transform -1 0 51520 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold135
timestamp 1704896540
transform -1 0 52256 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold136
timestamp 1704896540
transform 1 0 52716 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold137
timestamp 1704896540
transform 1 0 60352 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold138
timestamp 1704896540
transform -1 0 49680 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold139
timestamp 1704896540
transform -1 0 50784 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold140
timestamp 1704896540
transform 1 0 51152 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold141
timestamp 1704896540
transform 1 0 59340 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold142
timestamp 1704896540
transform 1 0 47104 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold143
timestamp 1704896540
transform -1 0 48944 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold144
timestamp 1704896540
transform 1 0 51336 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold145
timestamp 1704896540
transform -1 0 66332 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold146
timestamp 1704896540
transform 1 0 47104 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold147
timestamp 1704896540
transform 1 0 46368 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold148
timestamp 1704896540
transform 1 0 50600 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold149
timestamp 1704896540
transform -1 0 66332 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold150
timestamp 1704896540
transform -1 0 46368 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold151
timestamp 1704896540
transform 1 0 46000 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold152
timestamp 1704896540
transform 1 0 49864 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold153
timestamp 1704896540
transform -1 0 66332 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold154
timestamp 1704896540
transform 1 0 42320 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold155
timestamp 1704896540
transform -1 0 43792 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold156
timestamp 1704896540
transform 1 0 47564 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold157
timestamp 1704896540
transform -1 0 66332 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold158
timestamp 1704896540
transform -1 0 44528 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold159
timestamp 1704896540
transform -1 0 43056 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold160
timestamp 1704896540
transform 1 0 47840 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold161
timestamp 1704896540
transform -1 0 66332 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold162
timestamp 1704896540
transform 1 0 37444 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold163
timestamp 1704896540
transform -1 0 40480 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold164
timestamp 1704896540
transform 1 0 45448 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold165
timestamp 1704896540
transform -1 0 66332 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold166
timestamp 1704896540
transform -1 0 38548 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold167
timestamp 1704896540
transform -1 0 38732 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold168
timestamp 1704896540
transform 1 0 44252 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold169
timestamp 1704896540
transform -1 0 66332 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold170
timestamp 1704896540
transform 1 0 36156 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold171
timestamp 1704896540
transform 1 0 36248 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold172
timestamp 1704896540
transform 1 0 43424 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold173
timestamp 1704896540
transform -1 0 67804 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold174
timestamp 1704896540
transform -1 0 35788 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold175
timestamp 1704896540
transform 1 0 34684 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold176
timestamp 1704896540
transform 1 0 42228 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold177
timestamp 1704896540
transform -1 0 67068 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold178
timestamp 1704896540
transform 1 0 53360 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold179
timestamp 1704896540
transform -1 0 57408 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold180
timestamp 1704896540
transform -1 0 66332 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold181
timestamp 1704896540
transform -1 0 66332 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold182
timestamp 1704896540
transform -1 0 34316 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold183
timestamp 1704896540
transform -1 0 34040 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold184
timestamp 1704896540
transform 1 0 41308 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold185
timestamp 1704896540
transform -1 0 67804 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold186
timestamp 1704896540
transform 1 0 51612 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold187
timestamp 1704896540
transform -1 0 53084 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold188
timestamp 1704896540
transform 1 0 54372 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold189
timestamp 1704896540
transform -1 0 66332 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold190
timestamp 1704896540
transform 1 0 57776 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold191
timestamp 1704896540
transform -1 0 59984 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold192
timestamp 1704896540
transform -1 0 66332 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold193
timestamp 1704896540
transform -1 0 66332 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold194
timestamp 1704896540
transform 1 0 50784 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold195
timestamp 1704896540
transform -1 0 51888 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold196
timestamp 1704896540
transform 1 0 52992 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold197
timestamp 1704896540
transform -1 0 66332 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold198
timestamp 1704896540
transform -1 0 56672 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold199
timestamp 1704896540
transform -1 0 57408 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold200
timestamp 1704896540
transform -1 0 66332 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold201
timestamp 1704896540
transform -1 0 66332 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold202
timestamp 1704896540
transform 1 0 60352 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold203
timestamp 1704896540
transform -1 0 62560 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold204
timestamp 1704896540
transform -1 0 67068 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold205
timestamp 1704896540
transform -1 0 66332 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold206
timestamp 1704896540
transform 1 0 29256 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold207
timestamp 1704896540
transform -1 0 31096 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold208
timestamp 1704896540
transform 1 0 38548 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold209
timestamp 1704896540
transform -1 0 66332 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold210
timestamp 1704896540
transform 1 0 58880 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold211
timestamp 1704896540
transform 1 0 58512 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold212
timestamp 1704896540
transform -1 0 66332 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold213
timestamp 1704896540
transform -1 0 66332 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold214
timestamp 1704896540
transform 1 0 28612 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold215
timestamp 1704896540
transform 1 0 31188 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold216
timestamp 1704896540
transform 1 0 39928 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold217
timestamp 1704896540
transform -1 0 66332 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold218
timestamp 1704896540
transform 1 0 61088 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold219
timestamp 1704896540
transform -1 0 61456 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold220
timestamp 1704896540
transform 1 0 65596 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold221
timestamp 1704896540
transform -1 0 66332 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold222
timestamp 1704896540
transform 1 0 61456 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold223
timestamp 1704896540
transform -1 0 65136 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold224
timestamp 1704896540
transform 1 0 65596 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold225
timestamp 1704896540
transform -1 0 66332 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold226
timestamp 1704896540
transform -1 0 66240 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold227
timestamp 1704896540
transform -1 0 65136 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold228
timestamp 1704896540
transform -1 0 66332 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold229
timestamp 1704896540
transform -1 0 66332 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold230
timestamp 1704896540
transform -1 0 24196 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold231
timestamp 1704896540
transform 1 0 22724 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold232
timestamp 1704896540
transform 1 0 37168 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold233
timestamp 1704896540
transform -1 0 66332 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold234
timestamp 1704896540
transform 1 0 63112 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold235
timestamp 1704896540
transform 1 0 66792 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold236
timestamp 1704896540
transform 1 0 65596 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold237
timestamp 1704896540
transform -1 0 66332 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold238
timestamp 1704896540
transform 1 0 65596 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold239
timestamp 1704896540
transform 1 0 66976 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold240
timestamp 1704896540
transform -1 0 67068 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold241
timestamp 1704896540
transform -1 0 66332 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold242
timestamp 1704896540
transform -1 0 27600 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold243
timestamp 1704896540
transform -1 0 26036 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold244
timestamp 1704896540
transform 1 0 35696 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold245
timestamp 1704896540
transform -1 0 66332 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold246
timestamp 1704896540
transform -1 0 70288 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold247
timestamp 1704896540
transform 1 0 68448 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold248
timestamp 1704896540
transform -1 0 67804 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold249
timestamp 1704896540
transform -1 0 66332 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold250
timestamp 1704896540
transform -1 0 70840 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold251
timestamp 1704896540
transform -1 0 72864 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold252
timestamp 1704896540
transform -1 0 68908 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold253
timestamp 1704896540
transform -1 0 66332 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold254
timestamp 1704896540
transform 1 0 70656 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold255
timestamp 1704896540
transform -1 0 71116 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold256
timestamp 1704896540
transform -1 0 69368 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold257
timestamp 1704896540
transform -1 0 66332 0 -1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold258
timestamp 1704896540
transform 1 0 71208 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold259
timestamp 1704896540
transform -1 0 74704 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold260
timestamp 1704896540
transform -1 0 70840 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold261
timestamp 1704896540
transform -1 0 66424 0 1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold262
timestamp 1704896540
transform -1 0 45632 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold263
timestamp 1704896540
transform -1 0 46000 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold264
timestamp 1704896540
transform 1 0 48392 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold265
timestamp 1704896540
transform -1 0 67068 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold266
timestamp 1704896540
transform -1 0 42228 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold267
timestamp 1704896540
transform 1 0 43424 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold268
timestamp 1704896540
transform 1 0 47104 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold269
timestamp 1704896540
transform -1 0 66332 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold270
timestamp 1704896540
transform -1 0 41952 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold271
timestamp 1704896540
transform -1 0 41952 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold272
timestamp 1704896540
transform 1 0 46092 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold273
timestamp 1704896540
transform -1 0 67804 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold274
timestamp 1704896540
transform -1 0 39468 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold275
timestamp 1704896540
transform -1 0 39744 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold276
timestamp 1704896540
transform 1 0 44988 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold277
timestamp 1704896540
transform -1 0 67068 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold278
timestamp 1704896540
transform 1 0 35512 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold279
timestamp 1704896540
transform 1 0 37720 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold280
timestamp 1704896540
transform 1 0 44068 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold281
timestamp 1704896540
transform -1 0 67804 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold282
timestamp 1704896540
transform -1 0 35052 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold283
timestamp 1704896540
transform 1 0 33764 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold284
timestamp 1704896540
transform 1 0 41492 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold285
timestamp 1704896540
transform -1 0 66332 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold286
timestamp 1704896540
transform 1 0 34776 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold287
timestamp 1704896540
transform -1 0 36984 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold288
timestamp 1704896540
transform 1 0 42964 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold289
timestamp 1704896540
transform -1 0 66332 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold290
timestamp 1704896540
transform -1 0 30820 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold291
timestamp 1704896540
transform -1 0 33580 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold292
timestamp 1704896540
transform 1 0 40112 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold293
timestamp 1704896540
transform -1 0 66332 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold294
timestamp 1704896540
transform 1 0 28612 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold295
timestamp 1704896540
transform -1 0 30360 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold296
timestamp 1704896540
transform 1 0 38824 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold297
timestamp 1704896540
transform -1 0 66332 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold298
timestamp 1704896540
transform 1 0 25300 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold299
timestamp 1704896540
transform -1 0 29624 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold300
timestamp 1704896540
transform 1 0 38088 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold301
timestamp 1704896540
transform -1 0 66332 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold302
timestamp 1704896540
transform 1 0 21988 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold303
timestamp 1704896540
transform 1 0 26036 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold304
timestamp 1704896540
transform 1 0 26404 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold305
timestamp 1704896540
transform -1 0 25208 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold306
timestamp 1704896540
transform 1 0 23460 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold307
timestamp 1704896540
transform 1 0 32016 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold308
timestamp 1704896540
transform 1 0 35052 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold309
timestamp 1704896540
transform -1 0 28060 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold310
timestamp 1704896540
transform 1 0 22080 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold311
timestamp 1704896540
transform 1 0 20884 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold312
timestamp 1704896540
transform 1 0 24564 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold313
timestamp 1704896540
transform 1 0 49680 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold314
timestamp 1704896540
transform -1 0 50784 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold315
timestamp 1704896540
transform -1 0 52256 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold316
timestamp 1704896540
transform -1 0 49312 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold317
timestamp 1704896540
transform -1 0 48208 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold318
timestamp 1704896540
transform -1 0 50140 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold319
timestamp 1704896540
transform 1 0 45632 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold320
timestamp 1704896540
transform 1 0 47840 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold321
timestamp 1704896540
transform -1 0 46828 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold322
timestamp 1704896540
transform 1 0 44896 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold323
timestamp 1704896540
transform -1 0 44160 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold324
timestamp 1704896540
transform 1 0 43792 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold325
timestamp 1704896540
transform 1 0 41952 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold326
timestamp 1704896540
transform 1 0 41216 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold327
timestamp 1704896540
transform -1 0 41216 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold328
timestamp 1704896540
transform -1 0 41216 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold329
timestamp 1704896540
transform 1 0 36984 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold330
timestamp 1704896540
transform 1 0 36340 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold331
timestamp 1704896540
transform 1 0 34776 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold332
timestamp 1704896540
transform -1 0 37628 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold333
timestamp 1704896540
transform 1 0 34040 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold334
timestamp 1704896540
transform 1 0 32016 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold335
timestamp 1704896540
transform -1 0 55660 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold336
timestamp 1704896540
transform 1 0 54096 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold337
timestamp 1704896540
transform 1 0 29716 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold338
timestamp 1704896540
transform -1 0 33304 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold339
timestamp 1704896540
transform -1 0 53360 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold340
timestamp 1704896540
transform -1 0 54464 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold341
timestamp 1704896540
transform 1 0 54832 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold342
timestamp 1704896540
transform -1 0 55936 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold343
timestamp 1704896540
transform 1 0 56304 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold344
timestamp 1704896540
transform -1 0 58880 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold345
timestamp 1704896540
transform -1 0 54832 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold346
timestamp 1704896540
transform 1 0 52256 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold347
timestamp 1704896540
transform 1 0 57776 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold348
timestamp 1704896540
transform -1 0 61180 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold349
timestamp 1704896540
transform 1 0 59248 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold350
timestamp 1704896540
transform -1 0 30820 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold351
timestamp 1704896540
transform 1 0 59984 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold352
timestamp 1704896540
transform -1 0 30728 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold353
timestamp 1704896540
transform -1 0 62560 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold354
timestamp 1704896540
transform -1 0 64032 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold355
timestamp 1704896540
transform -1 0 25300 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold356
timestamp 1704896540
transform -1 0 66792 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold357
timestamp 1704896540
transform 1 0 25484 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold358
timestamp 1704896540
transform -1 0 66976 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold359
timestamp 1704896540
transform 1 0 67712 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold360
timestamp 1704896540
transform 1 0 69184 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold361
timestamp 1704896540
transform 1 0 69644 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold362
timestamp 1704896540
transform -1 0 73968 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold363
timestamp 1704896540
transform -1 0 47380 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold364
timestamp 1704896540
transform -1 0 43424 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold365
timestamp 1704896540
transform 1 0 40848 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold366
timestamp 1704896540
transform -1 0 41952 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold367
timestamp 1704896540
transform 1 0 34776 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold368
timestamp 1704896540
transform 1 0 32292 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold369
timestamp 1704896540
transform -1 0 36156 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold370
timestamp 1704896540
transform -1 0 32292 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold371
timestamp 1704896540
transform -1 0 26772 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold372
timestamp 1704896540
transform -1 0 31280 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1704896540
transform -1 0 21988 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input2
timestamp 1704896540
transform 1 0 44160 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input3
timestamp 1704896540
transform -1 0 44712 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input4
timestamp 1704896540
transform -1 0 29256 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input5
timestamp 1704896540
transform -1 0 28612 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input6
timestamp 1704896540
transform -1 0 30084 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input7
timestamp 1704896540
transform 1 0 34592 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input8
timestamp 1704896540
transform -1 0 36432 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input9
timestamp 1704896540
transform -1 0 37904 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input10
timestamp 1704896540
transform -1 0 39192 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input11
timestamp 1704896540
transform -1 0 40664 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1704896540
transform -1 0 24564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input13
timestamp 1704896540
transform -1 0 24932 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input14 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 42228 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input15 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 46828 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input16
timestamp 1704896540
transform 1 0 47472 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input17
timestamp 1704896540
transform -1 0 47104 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input18
timestamp 1704896540
transform -1 0 49680 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input19
timestamp 1704896540
transform -1 0 49680 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input20
timestamp 1704896540
transform -1 0 50692 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input21
timestamp 1704896540
transform -1 0 52440 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input22
timestamp 1704896540
transform -1 0 55016 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input23
timestamp 1704896540
transform -1 0 56212 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input24
timestamp 1704896540
transform 1 0 26864 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input25
timestamp 1704896540
transform -1 0 57592 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input26
timestamp 1704896540
transform -1 0 58788 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input27
timestamp 1704896540
transform -1 0 60168 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input28
timestamp 1704896540
transform -1 0 60996 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input29
timestamp 1704896540
transform -1 0 62744 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input30
timestamp 1704896540
transform 1 0 67344 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input31
timestamp 1704896540
transform -1 0 64584 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input32
timestamp 1704896540
transform 1 0 68080 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input33
timestamp 1704896540
transform -1 0 68632 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input34
timestamp 1704896540
transform -1 0 70472 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input35
timestamp 1704896540
transform -1 0 29992 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input36
timestamp 1704896540
transform 1 0 70840 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input37
timestamp 1704896540
transform -1 0 73784 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input38
timestamp 1704896540
transform 1 0 32016 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input39
timestamp 1704896540
transform -1 0 32568 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input40
timestamp 1704896540
transform 1 0 35144 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input41
timestamp 1704896540
transform -1 0 36984 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input42
timestamp 1704896540
transform -1 0 38180 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input43
timestamp 1704896540
transform -1 0 40020 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input44
timestamp 1704896540
transform -1 0 41216 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_12  input45
timestamp 1704896540
transform 1 0 27232 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  input46
timestamp 1704896540
transform 1 0 28980 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  input47
timestamp 1704896540
transform -1 0 31924 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  input48
timestamp 1704896540
transform 1 0 32752 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1704896540
transform -1 0 26036 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input50 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 26772 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__buf_12  output51
timestamp 1704896540
transform 1 0 24288 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output52
timestamp 1704896540
transform -1 0 28244 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output53
timestamp 1704896540
transform -1 0 43884 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output54
timestamp 1704896540
transform -1 0 45356 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output55
timestamp 1704896540
transform -1 0 46644 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output56
timestamp 1704896540
transform -1 0 48944 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output57
timestamp 1704896540
transform -1 0 49404 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output58
timestamp 1704896540
transform -1 0 51520 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output59
timestamp 1704896540
transform -1 0 52164 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output60
timestamp 1704896540
transform -1 0 54096 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output61
timestamp 1704896540
transform -1 0 54924 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output62
timestamp 1704896540
transform -1 0 56672 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output63
timestamp 1704896540
transform -1 0 29348 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output64
timestamp 1704896540
transform -1 0 57684 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output65
timestamp 1704896540
transform -1 0 59248 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output66
timestamp 1704896540
transform -1 0 60444 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output67
timestamp 1704896540
transform -1 0 61824 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output68
timestamp 1704896540
transform 1 0 62928 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output69
timestamp 1704896540
transform 1 0 63112 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output70
timestamp 1704896540
transform 1 0 64584 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output71
timestamp 1704896540
transform 1 0 65872 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output72
timestamp 1704896540
transform 1 0 68080 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output73
timestamp 1704896540
transform 1 0 68632 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output74
timestamp 1704896540
transform -1 0 31924 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output75
timestamp 1704896540
transform 1 0 70656 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output76
timestamp 1704896540
transform 1 0 71392 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output77
timestamp 1704896540
transform -1 0 33764 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output78
timestamp 1704896540
transform -1 0 35604 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output79
timestamp 1704896540
transform -1 0 36984 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output80
timestamp 1704896540
transform -1 0 38640 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output81
timestamp 1704896540
transform -1 0 39652 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output82
timestamp 1704896540
transform -1 0 41216 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output83
timestamp 1704896540
transform -1 0 43792 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_0
timestamp 1704896540
transform 1 0 1012 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_9
timestamp 1704896540
transform -1 0 74980 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_1
timestamp 1704896540
transform 1 0 1012 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_10
timestamp 1704896540
transform -1 0 74980 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_2
timestamp 1704896540
transform 1 0 1012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_11
timestamp 1704896540
transform -1 0 74980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_3
timestamp 1704896540
transform 1 0 1012 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_12
timestamp 1704896540
transform -1 0 74980 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_4
timestamp 1704896540
transform 1 0 1012 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_13
timestamp 1704896540
transform -1 0 74980 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_5
timestamp 1704896540
transform 1 0 1012 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_14
timestamp 1704896540
transform -1 0 74980 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_6
timestamp 1704896540
transform 1 0 1012 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_15
timestamp 1704896540
transform -1 0 74980 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_7
timestamp 1704896540
transform 1 0 1012 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_16
timestamp 1704896540
transform -1 0 74980 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_8
timestamp 1704896540
transform 1 0 1012 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_17
timestamp 1704896540
transform -1 0 74980 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_2_Left_311
timestamp 1704896540
transform 1 0 65320 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_2_Right_164
timestamp 1704896540
transform -1 0 74980 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_2_Left_165
timestamp 1704896540
transform 1 0 65320 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_2_Right_18
timestamp 1704896540
transform -1 0 74980 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_2_Left_166
timestamp 1704896540
transform 1 0 65320 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_2_Right_19
timestamp 1704896540
transform -1 0 74980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_2_Left_167
timestamp 1704896540
transform 1 0 65320 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_2_Right_20
timestamp 1704896540
transform -1 0 74980 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_2_Left_168
timestamp 1704896540
transform 1 0 65320 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_2_Right_21
timestamp 1704896540
transform -1 0 74980 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_2_Left_169
timestamp 1704896540
transform 1 0 65320 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_2_Right_22
timestamp 1704896540
transform -1 0 74980 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_2_Left_170
timestamp 1704896540
transform 1 0 65320 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_2_Right_23
timestamp 1704896540
transform -1 0 74980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_2_Left_171
timestamp 1704896540
transform 1 0 65320 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_2_Right_24
timestamp 1704896540
transform -1 0 74980 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_2_Left_172
timestamp 1704896540
transform 1 0 65320 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_2_Right_25
timestamp 1704896540
transform -1 0 74980 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_2_Left_173
timestamp 1704896540
transform 1 0 65320 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_2_Right_26
timestamp 1704896540
transform -1 0 74980 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_2_Left_174
timestamp 1704896540
transform 1 0 65320 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_2_Right_27
timestamp 1704896540
transform -1 0 74980 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_2_Left_175
timestamp 1704896540
transform 1 0 65320 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_2_Right_28
timestamp 1704896540
transform -1 0 74980 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_2_Left_176
timestamp 1704896540
transform 1 0 65320 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_2_Right_29
timestamp 1704896540
transform -1 0 74980 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_2_Left_177
timestamp 1704896540
transform 1 0 65320 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_2_Right_30
timestamp 1704896540
transform -1 0 74980 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_2_Left_178
timestamp 1704896540
transform 1 0 65320 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_2_Right_31
timestamp 1704896540
transform -1 0 74980 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_2_Left_179
timestamp 1704896540
transform 1 0 65320 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_2_Right_32
timestamp 1704896540
transform -1 0 74980 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_2_Left_180
timestamp 1704896540
transform 1 0 65320 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_2_Right_33
timestamp 1704896540
transform -1 0 74980 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_2_Left_181
timestamp 1704896540
transform 1 0 65320 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_2_Right_34
timestamp 1704896540
transform -1 0 74980 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_2_Left_182
timestamp 1704896540
transform 1 0 65320 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_2_Right_35
timestamp 1704896540
transform -1 0 74980 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_2_Left_183
timestamp 1704896540
transform 1 0 65320 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_2_Right_36
timestamp 1704896540
transform -1 0 74980 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_2_Left_184
timestamp 1704896540
transform 1 0 65320 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_2_Right_37
timestamp 1704896540
transform -1 0 74980 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_2_Left_185
timestamp 1704896540
transform 1 0 65320 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_2_Right_38
timestamp 1704896540
transform -1 0 74980 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_2_Left_186
timestamp 1704896540
transform 1 0 65320 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_2_Right_39
timestamp 1704896540
transform -1 0 74980 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_2_Left_187
timestamp 1704896540
transform 1 0 65320 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_2_Right_40
timestamp 1704896540
transform -1 0 74980 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_2_Left_188
timestamp 1704896540
transform 1 0 65320 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_2_Right_41
timestamp 1704896540
transform -1 0 74980 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_2_Left_189
timestamp 1704896540
transform 1 0 65320 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_2_Right_42
timestamp 1704896540
transform -1 0 74980 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_2_Left_190
timestamp 1704896540
transform 1 0 65320 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_2_Right_43
timestamp 1704896540
transform -1 0 74980 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_2_Left_191
timestamp 1704896540
transform 1 0 65320 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_2_Right_44
timestamp 1704896540
transform -1 0 74980 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_2_Left_192
timestamp 1704896540
transform 1 0 65320 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_2_Right_45
timestamp 1704896540
transform -1 0 74980 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_2_Left_193
timestamp 1704896540
transform 1 0 65320 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_2_Right_46
timestamp 1704896540
transform -1 0 74980 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_2_Left_194
timestamp 1704896540
transform 1 0 65320 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_2_Right_47
timestamp 1704896540
transform -1 0 74980 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_2_Left_195
timestamp 1704896540
transform 1 0 65320 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_2_Right_48
timestamp 1704896540
transform -1 0 74980 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_2_Left_196
timestamp 1704896540
transform 1 0 65320 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_2_Right_49
timestamp 1704896540
transform -1 0 74980 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_2_Left_197
timestamp 1704896540
transform 1 0 65320 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_2_Right_50
timestamp 1704896540
transform -1 0 74980 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_2_Left_198
timestamp 1704896540
transform 1 0 65320 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_2_Right_51
timestamp 1704896540
transform -1 0 74980 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_2_Left_199
timestamp 1704896540
transform 1 0 65320 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_2_Right_52
timestamp 1704896540
transform -1 0 74980 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_2_Left_200
timestamp 1704896540
transform 1 0 65320 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_2_Right_53
timestamp 1704896540
transform -1 0 74980 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_2_Left_201
timestamp 1704896540
transform 1 0 65320 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_2_Right_54
timestamp 1704896540
transform -1 0 74980 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_2_Left_202
timestamp 1704896540
transform 1 0 65320 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_2_Right_55
timestamp 1704896540
transform -1 0 74980 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_2_Left_203
timestamp 1704896540
transform 1 0 65320 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_2_Right_56
timestamp 1704896540
transform -1 0 74980 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_2_Left_204
timestamp 1704896540
transform 1 0 65320 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_2_Right_57
timestamp 1704896540
transform -1 0 74980 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_2_Left_205
timestamp 1704896540
transform 1 0 65320 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_2_Right_58
timestamp 1704896540
transform -1 0 74980 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_2_Left_206
timestamp 1704896540
transform 1 0 65320 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_2_Right_59
timestamp 1704896540
transform -1 0 74980 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_2_Left_207
timestamp 1704896540
transform 1 0 65320 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_2_Right_60
timestamp 1704896540
transform -1 0 74980 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_2_Left_208
timestamp 1704896540
transform 1 0 65320 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_2_Right_61
timestamp 1704896540
transform -1 0 74980 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_2_Left_209
timestamp 1704896540
transform 1 0 65320 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_2_Right_62
timestamp 1704896540
transform -1 0 74980 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_2_Left_210
timestamp 1704896540
transform 1 0 65320 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_2_Right_63
timestamp 1704896540
transform -1 0 74980 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_2_Left_211
timestamp 1704896540
transform 1 0 65320 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_2_Right_64
timestamp 1704896540
transform -1 0 74980 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_2_Left_212
timestamp 1704896540
transform 1 0 65320 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_2_Right_65
timestamp 1704896540
transform -1 0 74980 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_2_Left_213
timestamp 1704896540
transform 1 0 65320 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_2_Right_66
timestamp 1704896540
transform -1 0 74980 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_2_Left_214
timestamp 1704896540
transform 1 0 65320 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_2_Right_67
timestamp 1704896540
transform -1 0 74980 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_2_Left_215
timestamp 1704896540
transform 1 0 65320 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_2_Right_68
timestamp 1704896540
transform -1 0 74980 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_2_Left_216
timestamp 1704896540
transform 1 0 65320 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_2_Right_69
timestamp 1704896540
transform -1 0 74980 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_2_Left_217
timestamp 1704896540
transform 1 0 65320 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_2_Right_70
timestamp 1704896540
transform -1 0 74980 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_2_Left_218
timestamp 1704896540
transform 1 0 65320 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_2_Right_71
timestamp 1704896540
transform -1 0 74980 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_2_Left_219
timestamp 1704896540
transform 1 0 65320 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_2_Right_72
timestamp 1704896540
transform -1 0 74980 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_2_Left_220
timestamp 1704896540
transform 1 0 65320 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_2_Right_73
timestamp 1704896540
transform -1 0 74980 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_2_Left_221
timestamp 1704896540
transform 1 0 65320 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_2_Right_74
timestamp 1704896540
transform -1 0 74980 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_2_Left_222
timestamp 1704896540
transform 1 0 65320 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_2_Right_75
timestamp 1704896540
transform -1 0 74980 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_2_Left_223
timestamp 1704896540
transform 1 0 65320 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_2_Right_76
timestamp 1704896540
transform -1 0 74980 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_2_Left_224
timestamp 1704896540
transform 1 0 65320 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_2_Right_77
timestamp 1704896540
transform -1 0 74980 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_2_Left_225
timestamp 1704896540
transform 1 0 65320 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_2_Right_78
timestamp 1704896540
transform -1 0 74980 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_2_Left_226
timestamp 1704896540
transform 1 0 65320 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_2_Right_79
timestamp 1704896540
transform -1 0 74980 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_2_Left_227
timestamp 1704896540
transform 1 0 65320 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_2_Right_80
timestamp 1704896540
transform -1 0 74980 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_2_Left_228
timestamp 1704896540
transform 1 0 65320 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_2_Right_81
timestamp 1704896540
transform -1 0 74980 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_2_Left_229
timestamp 1704896540
transform 1 0 65320 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_2_Right_82
timestamp 1704896540
transform -1 0 74980 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_2_Left_230
timestamp 1704896540
transform 1 0 65320 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_2_Right_83
timestamp 1704896540
transform -1 0 74980 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_2_Left_231
timestamp 1704896540
transform 1 0 65320 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_2_Right_84
timestamp 1704896540
transform -1 0 74980 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_2_Left_232
timestamp 1704896540
transform 1 0 65320 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_2_Right_85
timestamp 1704896540
transform -1 0 74980 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_2_Left_233
timestamp 1704896540
transform 1 0 65320 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_2_Right_86
timestamp 1704896540
transform -1 0 74980 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_2_Left_234
timestamp 1704896540
transform 1 0 65320 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_2_Right_87
timestamp 1704896540
transform -1 0 74980 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_2_Left_235
timestamp 1704896540
transform 1 0 65320 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_2_Right_88
timestamp 1704896540
transform -1 0 74980 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_2_Left_236
timestamp 1704896540
transform 1 0 65320 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_2_Right_89
timestamp 1704896540
transform -1 0 74980 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_2_Left_237
timestamp 1704896540
transform 1 0 65320 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_2_Right_90
timestamp 1704896540
transform -1 0 74980 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_2_Left_238
timestamp 1704896540
transform 1 0 65320 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_2_Right_91
timestamp 1704896540
transform -1 0 74980 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_2_Left_239
timestamp 1704896540
transform 1 0 65320 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_2_Right_92
timestamp 1704896540
transform -1 0 74980 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_2_Left_240
timestamp 1704896540
transform 1 0 65320 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_2_Right_93
timestamp 1704896540
transform -1 0 74980 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_2_Left_241
timestamp 1704896540
transform 1 0 65320 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_2_Right_94
timestamp 1704896540
transform -1 0 74980 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_2_Left_242
timestamp 1704896540
transform 1 0 65320 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_2_Right_95
timestamp 1704896540
transform -1 0 74980 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_2_Left_243
timestamp 1704896540
transform 1 0 65320 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_2_Right_96
timestamp 1704896540
transform -1 0 74980 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_2_Left_244
timestamp 1704896540
transform 1 0 65320 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_2_Right_97
timestamp 1704896540
transform -1 0 74980 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_2_Left_245
timestamp 1704896540
transform 1 0 65320 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_2_Right_98
timestamp 1704896540
transform -1 0 74980 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_2_Left_246
timestamp 1704896540
transform 1 0 65320 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_2_Right_99
timestamp 1704896540
transform -1 0 74980 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_2_Left_247
timestamp 1704896540
transform 1 0 65320 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_2_Right_100
timestamp 1704896540
transform -1 0 74980 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_2_Left_248
timestamp 1704896540
transform 1 0 65320 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_2_Right_101
timestamp 1704896540
transform -1 0 74980 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_2_Left_249
timestamp 1704896540
transform 1 0 65320 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_2_Right_102
timestamp 1704896540
transform -1 0 74980 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_2_Left_250
timestamp 1704896540
transform 1 0 65320 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_2_Right_103
timestamp 1704896540
transform -1 0 74980 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_2_Left_251
timestamp 1704896540
transform 1 0 65320 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_2_Right_104
timestamp 1704896540
transform -1 0 74980 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_2_Left_252
timestamp 1704896540
transform 1 0 65320 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_2_Right_105
timestamp 1704896540
transform -1 0 74980 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_2_Left_253
timestamp 1704896540
transform 1 0 65320 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_2_Right_106
timestamp 1704896540
transform -1 0 74980 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_2_Left_254
timestamp 1704896540
transform 1 0 65320 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_2_Right_107
timestamp 1704896540
transform -1 0 74980 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_2_Left_255
timestamp 1704896540
transform 1 0 65320 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_2_Right_108
timestamp 1704896540
transform -1 0 74980 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_2_Left_256
timestamp 1704896540
transform 1 0 65320 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_2_Right_109
timestamp 1704896540
transform -1 0 74980 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_2_Left_257
timestamp 1704896540
transform 1 0 65320 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_2_Right_110
timestamp 1704896540
transform -1 0 74980 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_2_Left_258
timestamp 1704896540
transform 1 0 65320 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_2_Right_111
timestamp 1704896540
transform -1 0 74980 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_2_Left_259
timestamp 1704896540
transform 1 0 65320 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_2_Right_112
timestamp 1704896540
transform -1 0 74980 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_2_Left_260
timestamp 1704896540
transform 1 0 65320 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_2_Right_113
timestamp 1704896540
transform -1 0 74980 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_2_Left_261
timestamp 1704896540
transform 1 0 65320 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_2_Right_114
timestamp 1704896540
transform -1 0 74980 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_2_Left_262
timestamp 1704896540
transform 1 0 65320 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_2_Right_115
timestamp 1704896540
transform -1 0 74980 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_2_Left_263
timestamp 1704896540
transform 1 0 65320 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_2_Right_116
timestamp 1704896540
transform -1 0 74980 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_2_Left_264
timestamp 1704896540
transform 1 0 65320 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_2_Right_117
timestamp 1704896540
transform -1 0 74980 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_2_Left_265
timestamp 1704896540
transform 1 0 65320 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_2_Right_118
timestamp 1704896540
transform -1 0 74980 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_2_Left_266
timestamp 1704896540
transform 1 0 65320 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_2_Right_119
timestamp 1704896540
transform -1 0 74980 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_2_Left_267
timestamp 1704896540
transform 1 0 65320 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_2_Right_120
timestamp 1704896540
transform -1 0 74980 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_2_Left_268
timestamp 1704896540
transform 1 0 65320 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_2_Right_121
timestamp 1704896540
transform -1 0 74980 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_2_Left_269
timestamp 1704896540
transform 1 0 65320 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_2_Right_122
timestamp 1704896540
transform -1 0 74980 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_2_Left_270
timestamp 1704896540
transform 1 0 65320 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_2_Right_123
timestamp 1704896540
transform -1 0 74980 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_2_Left_271
timestamp 1704896540
transform 1 0 65320 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_2_Right_124
timestamp 1704896540
transform -1 0 74980 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_117_2_Left_272
timestamp 1704896540
transform 1 0 65320 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_117_2_Right_125
timestamp 1704896540
transform -1 0 74980 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_118_2_Left_273
timestamp 1704896540
transform 1 0 65320 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_118_2_Right_126
timestamp 1704896540
transform -1 0 74980 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_119_2_Left_274
timestamp 1704896540
transform 1 0 65320 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_119_2_Right_127
timestamp 1704896540
transform -1 0 74980 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_120_2_Left_275
timestamp 1704896540
transform 1 0 65320 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_120_2_Right_128
timestamp 1704896540
transform -1 0 74980 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_2_Left_276
timestamp 1704896540
transform 1 0 65320 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_2_Right_129
timestamp 1704896540
transform -1 0 74980 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_2_Left_277
timestamp 1704896540
transform 1 0 65320 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_2_Right_130
timestamp 1704896540
transform -1 0 74980 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_2_Left_278
timestamp 1704896540
transform 1 0 65320 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_2_Right_131
timestamp 1704896540
transform -1 0 74980 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_124_2_Left_279
timestamp 1704896540
transform 1 0 65320 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_124_2_Right_132
timestamp 1704896540
transform -1 0 74980 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_125_2_Left_280
timestamp 1704896540
transform 1 0 65320 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_125_2_Right_133
timestamp 1704896540
transform -1 0 74980 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_126_2_Left_281
timestamp 1704896540
transform 1 0 65320 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_126_2_Right_134
timestamp 1704896540
transform -1 0 74980 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_127_2_Left_282
timestamp 1704896540
transform 1 0 65320 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_127_2_Right_135
timestamp 1704896540
transform -1 0 74980 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_128_2_Left_283
timestamp 1704896540
transform 1 0 65320 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_128_2_Right_136
timestamp 1704896540
transform -1 0 74980 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_129_2_Left_284
timestamp 1704896540
transform 1 0 65320 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_129_2_Right_137
timestamp 1704896540
transform -1 0 74980 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_130_2_Left_285
timestamp 1704896540
transform 1 0 65320 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_130_2_Right_138
timestamp 1704896540
transform -1 0 74980 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_131_2_Left_286
timestamp 1704896540
transform 1 0 65320 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_131_2_Right_139
timestamp 1704896540
transform -1 0 74980 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_132_2_Left_287
timestamp 1704896540
transform 1 0 65320 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_132_2_Right_140
timestamp 1704896540
transform -1 0 74980 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_133_2_Left_288
timestamp 1704896540
transform 1 0 65320 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_133_2_Right_141
timestamp 1704896540
transform -1 0 74980 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_134_2_Left_289
timestamp 1704896540
transform 1 0 65320 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_134_2_Right_142
timestamp 1704896540
transform -1 0 74980 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_135_2_Left_290
timestamp 1704896540
transform 1 0 65320 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_135_2_Right_143
timestamp 1704896540
transform -1 0 74980 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_136_2_Left_291
timestamp 1704896540
transform 1 0 65320 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_136_2_Right_144
timestamp 1704896540
transform -1 0 74980 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_137_2_Left_292
timestamp 1704896540
transform 1 0 65320 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_137_2_Right_145
timestamp 1704896540
transform -1 0 74980 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_138_2_Left_293
timestamp 1704896540
transform 1 0 65320 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_138_2_Right_146
timestamp 1704896540
transform -1 0 74980 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_139_2_Left_294
timestamp 1704896540
transform 1 0 65320 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_139_2_Right_147
timestamp 1704896540
transform -1 0 74980 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_140_2_Left_295
timestamp 1704896540
transform 1 0 65320 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_140_2_Right_148
timestamp 1704896540
transform -1 0 74980 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_141_2_Left_296
timestamp 1704896540
transform 1 0 65320 0 -1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_141_2_Right_149
timestamp 1704896540
transform -1 0 74980 0 -1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_142_2_Left_297
timestamp 1704896540
transform 1 0 65320 0 1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_142_2_Right_150
timestamp 1704896540
transform -1 0 74980 0 1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_143_2_Left_298
timestamp 1704896540
transform 1 0 65320 0 -1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_143_2_Right_151
timestamp 1704896540
transform -1 0 74980 0 -1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_144_2_Left_299
timestamp 1704896540
transform 1 0 65320 0 1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_144_2_Right_152
timestamp 1704896540
transform -1 0 74980 0 1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_145_2_Left_300
timestamp 1704896540
transform 1 0 65320 0 -1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_145_2_Right_153
timestamp 1704896540
transform -1 0 74980 0 -1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_146_2_Left_301
timestamp 1704896540
transform 1 0 65320 0 1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_146_2_Right_154
timestamp 1704896540
transform -1 0 74980 0 1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_147_2_Left_302
timestamp 1704896540
transform 1 0 65320 0 -1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_147_2_Right_155
timestamp 1704896540
transform -1 0 74980 0 -1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_148_2_Left_303
timestamp 1704896540
transform 1 0 65320 0 1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_148_2_Right_156
timestamp 1704896540
transform -1 0 74980 0 1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_149_2_Left_304
timestamp 1704896540
transform 1 0 65320 0 -1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_149_2_Right_157
timestamp 1704896540
transform -1 0 74980 0 -1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_150_2_Left_305
timestamp 1704896540
transform 1 0 65320 0 1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_150_2_Right_158
timestamp 1704896540
transform -1 0 74980 0 1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_151_2_Left_306
timestamp 1704896540
transform 1 0 65320 0 -1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_151_2_Right_159
timestamp 1704896540
transform -1 0 74980 0 -1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_152_2_Left_307
timestamp 1704896540
transform 1 0 65320 0 1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_152_2_Right_160
timestamp 1704896540
transform -1 0 74980 0 1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_153_2_Left_308
timestamp 1704896540
transform 1 0 65320 0 -1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_153_2_Right_161
timestamp 1704896540
transform -1 0 74980 0 -1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_154_2_Left_309
timestamp 1704896540
transform 1 0 65320 0 1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_154_2_Right_162
timestamp 1704896540
transform -1 0 74980 0 1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_155_2_Left_310
timestamp 1704896540
transform 1 0 65320 0 -1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_155_2_Right_163
timestamp 1704896540
transform -1 0 74980 0 -1 85952
box -38 -48 314 592
use EF_SRAM_1024x32  SRAM_0
timestamp 0
transform 0 -1 63283 1 0 8000
box 0 -40 77574 61263
use sky130_fd_sc_hd__conb_1  SRAM_0_84 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 65872 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  SRAM_0_85
timestamp 1704896540
transform -1 0 66608 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  SRAM_0_86
timestamp 1704896540
transform -1 0 65872 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  SRAM_0_87
timestamp 1704896540
transform -1 0 66608 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  SRAM_0_88
timestamp 1704896540
transform -1 0 65872 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  SRAM_0_89
timestamp 1704896540
transform -1 0 66148 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  SRAM_0_90
timestamp 1704896540
transform -1 0 65872 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  SRAM_0_91
timestamp 1704896540
transform 1 0 66332 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  SRAM_0_92
timestamp 1704896540
transform 1 0 66608 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_312 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3588 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_313
timestamp 1704896540
transform 1 0 6164 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_314
timestamp 1704896540
transform 1 0 8740 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_315
timestamp 1704896540
transform 1 0 11316 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_316
timestamp 1704896540
transform 1 0 13892 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_317
timestamp 1704896540
transform 1 0 16468 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_318
timestamp 1704896540
transform 1 0 19044 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_319
timestamp 1704896540
transform 1 0 21620 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_320
timestamp 1704896540
transform 1 0 24196 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_321
timestamp 1704896540
transform 1 0 26772 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_322
timestamp 1704896540
transform 1 0 29348 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_323
timestamp 1704896540
transform 1 0 31924 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_324
timestamp 1704896540
transform 1 0 34500 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_325
timestamp 1704896540
transform 1 0 37076 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_326
timestamp 1704896540
transform 1 0 39652 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_327
timestamp 1704896540
transform 1 0 42228 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_328
timestamp 1704896540
transform 1 0 44804 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_329
timestamp 1704896540
transform 1 0 47380 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_330
timestamp 1704896540
transform 1 0 49956 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_331
timestamp 1704896540
transform 1 0 52532 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_332
timestamp 1704896540
transform 1 0 55108 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_333
timestamp 1704896540
transform 1 0 57684 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_334
timestamp 1704896540
transform 1 0 60260 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_335
timestamp 1704896540
transform 1 0 62836 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_336
timestamp 1704896540
transform 1 0 65412 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_337
timestamp 1704896540
transform 1 0 67988 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_338
timestamp 1704896540
transform 1 0 70564 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_339
timestamp 1704896540
transform 1 0 73140 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_340
timestamp 1704896540
transform 1 0 6164 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_341
timestamp 1704896540
transform 1 0 11316 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_342
timestamp 1704896540
transform 1 0 16468 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_343
timestamp 1704896540
transform 1 0 21620 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_344
timestamp 1704896540
transform 1 0 26772 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_345
timestamp 1704896540
transform 1 0 31924 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_346
timestamp 1704896540
transform 1 0 37076 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_347
timestamp 1704896540
transform 1 0 42228 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_348
timestamp 1704896540
transform 1 0 47380 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_349
timestamp 1704896540
transform 1 0 52532 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_350
timestamp 1704896540
transform 1 0 57684 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_351
timestamp 1704896540
transform 1 0 62836 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_352
timestamp 1704896540
transform 1 0 67988 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_353
timestamp 1704896540
transform 1 0 73140 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_354
timestamp 1704896540
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_355
timestamp 1704896540
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_356
timestamp 1704896540
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_357
timestamp 1704896540
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_358
timestamp 1704896540
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_359
timestamp 1704896540
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_360
timestamp 1704896540
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_361
timestamp 1704896540
transform 1 0 39652 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_362
timestamp 1704896540
transform 1 0 44804 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_363
timestamp 1704896540
transform 1 0 49956 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_364
timestamp 1704896540
transform 1 0 55108 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_365
timestamp 1704896540
transform 1 0 60260 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_366
timestamp 1704896540
transform 1 0 65412 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_367
timestamp 1704896540
transform 1 0 70564 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_368
timestamp 1704896540
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_369
timestamp 1704896540
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_370
timestamp 1704896540
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_371
timestamp 1704896540
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_372
timestamp 1704896540
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_373
timestamp 1704896540
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_374
timestamp 1704896540
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_375
timestamp 1704896540
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_376
timestamp 1704896540
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_377
timestamp 1704896540
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_378
timestamp 1704896540
transform 1 0 57684 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_379
timestamp 1704896540
transform 1 0 62836 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_380
timestamp 1704896540
transform 1 0 67988 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_381
timestamp 1704896540
transform 1 0 73140 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_382
timestamp 1704896540
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_383
timestamp 1704896540
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_384
timestamp 1704896540
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_385
timestamp 1704896540
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_386
timestamp 1704896540
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_387
timestamp 1704896540
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_388
timestamp 1704896540
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_389
timestamp 1704896540
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_390
timestamp 1704896540
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_391
timestamp 1704896540
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_392
timestamp 1704896540
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_393
timestamp 1704896540
transform 1 0 60260 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_394
timestamp 1704896540
transform 1 0 65412 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_395
timestamp 1704896540
transform 1 0 70564 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_396
timestamp 1704896540
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_397
timestamp 1704896540
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_398
timestamp 1704896540
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_399
timestamp 1704896540
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_400
timestamp 1704896540
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_401
timestamp 1704896540
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_402
timestamp 1704896540
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_403
timestamp 1704896540
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_404
timestamp 1704896540
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_405
timestamp 1704896540
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_406
timestamp 1704896540
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_407
timestamp 1704896540
transform 1 0 62836 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_408
timestamp 1704896540
transform 1 0 67988 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_409
timestamp 1704896540
transform 1 0 73140 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_410
timestamp 1704896540
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_411
timestamp 1704896540
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_412
timestamp 1704896540
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_413
timestamp 1704896540
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_414
timestamp 1704896540
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_415
timestamp 1704896540
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_416
timestamp 1704896540
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_417
timestamp 1704896540
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_418
timestamp 1704896540
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_419
timestamp 1704896540
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_420
timestamp 1704896540
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_421
timestamp 1704896540
transform 1 0 60260 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_422
timestamp 1704896540
transform 1 0 65412 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_423
timestamp 1704896540
transform 1 0 70564 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_424
timestamp 1704896540
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_425
timestamp 1704896540
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_426
timestamp 1704896540
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_427
timestamp 1704896540
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_428
timestamp 1704896540
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_429
timestamp 1704896540
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_430
timestamp 1704896540
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_431
timestamp 1704896540
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_432
timestamp 1704896540
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_433
timestamp 1704896540
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_434
timestamp 1704896540
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_435
timestamp 1704896540
transform 1 0 62836 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_436
timestamp 1704896540
transform 1 0 67988 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_437
timestamp 1704896540
transform 1 0 73140 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_438
timestamp 1704896540
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_439
timestamp 1704896540
transform 1 0 6164 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_440
timestamp 1704896540
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_441
timestamp 1704896540
transform 1 0 11316 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_442
timestamp 1704896540
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_443
timestamp 1704896540
transform 1 0 16468 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_444
timestamp 1704896540
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_445
timestamp 1704896540
transform 1 0 21620 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_446
timestamp 1704896540
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_447
timestamp 1704896540
transform 1 0 26772 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_448
timestamp 1704896540
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_449
timestamp 1704896540
transform 1 0 31924 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_450
timestamp 1704896540
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_451
timestamp 1704896540
transform 1 0 37076 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_452
timestamp 1704896540
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_453
timestamp 1704896540
transform 1 0 42228 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_454
timestamp 1704896540
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_455
timestamp 1704896540
transform 1 0 47380 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_456
timestamp 1704896540
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_457
timestamp 1704896540
transform 1 0 52532 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_458
timestamp 1704896540
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_459
timestamp 1704896540
transform 1 0 57684 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_460
timestamp 1704896540
transform 1 0 60260 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_461
timestamp 1704896540
transform 1 0 62836 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_462
timestamp 1704896540
transform 1 0 65412 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_463
timestamp 1704896540
transform 1 0 67988 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_464
timestamp 1704896540
transform 1 0 70564 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_465
timestamp 1704896540
transform 1 0 73140 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_2_687
timestamp 1704896540
transform 1 0 70472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_2_466
timestamp 1704896540
transform 1 0 67896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_2_467
timestamp 1704896540
transform 1 0 73048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_2_468
timestamp 1704896540
transform 1 0 70472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_2_469
timestamp 1704896540
transform 1 0 67896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_2_470
timestamp 1704896540
transform 1 0 73048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_2_471
timestamp 1704896540
transform 1 0 70472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_2_472
timestamp 1704896540
transform 1 0 67896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_2_473
timestamp 1704896540
transform 1 0 73048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_2_474
timestamp 1704896540
transform 1 0 70472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_2_475
timestamp 1704896540
transform 1 0 67896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_2_476
timestamp 1704896540
transform 1 0 73048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_2_477
timestamp 1704896540
transform 1 0 70472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_2_478
timestamp 1704896540
transform 1 0 67896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_2_479
timestamp 1704896540
transform 1 0 73048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_2_480
timestamp 1704896540
transform 1 0 70472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_2_481
timestamp 1704896540
transform 1 0 67896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_2_482
timestamp 1704896540
transform 1 0 73048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_2_483
timestamp 1704896540
transform 1 0 70472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_2_484
timestamp 1704896540
transform 1 0 67896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_2_485
timestamp 1704896540
transform 1 0 73048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_2_486
timestamp 1704896540
transform 1 0 70472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_2_487
timestamp 1704896540
transform 1 0 67896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_2_488
timestamp 1704896540
transform 1 0 73048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_2_489
timestamp 1704896540
transform 1 0 70472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_2_490
timestamp 1704896540
transform 1 0 67896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_2_491
timestamp 1704896540
transform 1 0 73048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_2_492
timestamp 1704896540
transform 1 0 70472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_2_493
timestamp 1704896540
transform 1 0 67896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_2_494
timestamp 1704896540
transform 1 0 73048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_2_495
timestamp 1704896540
transform 1 0 70472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_2_496
timestamp 1704896540
transform 1 0 67896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_2_497
timestamp 1704896540
transform 1 0 73048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_2_498
timestamp 1704896540
transform 1 0 70472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_2_499
timestamp 1704896540
transform 1 0 67896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_2_500
timestamp 1704896540
transform 1 0 73048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_2_501
timestamp 1704896540
transform 1 0 70472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_2_502
timestamp 1704896540
transform 1 0 67896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_2_503
timestamp 1704896540
transform 1 0 73048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_2_504
timestamp 1704896540
transform 1 0 70472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_2_505
timestamp 1704896540
transform 1 0 67896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_2_506
timestamp 1704896540
transform 1 0 73048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_2_507
timestamp 1704896540
transform 1 0 70472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_2_508
timestamp 1704896540
transform 1 0 67896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_2_509
timestamp 1704896540
transform 1 0 73048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_2_510
timestamp 1704896540
transform 1 0 70472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_2_511
timestamp 1704896540
transform 1 0 67896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_2_512
timestamp 1704896540
transform 1 0 73048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_2_513
timestamp 1704896540
transform 1 0 70472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_2_514
timestamp 1704896540
transform 1 0 67896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_2_515
timestamp 1704896540
transform 1 0 73048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_2_516
timestamp 1704896540
transform 1 0 70472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_2_517
timestamp 1704896540
transform 1 0 67896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_2_518
timestamp 1704896540
transform 1 0 73048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_2_519
timestamp 1704896540
transform 1 0 70472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_2_520
timestamp 1704896540
transform 1 0 67896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_2_521
timestamp 1704896540
transform 1 0 73048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_2_522
timestamp 1704896540
transform 1 0 70472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_2_523
timestamp 1704896540
transform 1 0 67896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_2_524
timestamp 1704896540
transform 1 0 73048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_2_525
timestamp 1704896540
transform 1 0 70472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_2_526
timestamp 1704896540
transform 1 0 67896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_2_527
timestamp 1704896540
transform 1 0 73048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_2_528
timestamp 1704896540
transform 1 0 70472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_2_529
timestamp 1704896540
transform 1 0 67896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_2_530
timestamp 1704896540
transform 1 0 73048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_2_531
timestamp 1704896540
transform 1 0 70472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_2_532
timestamp 1704896540
transform 1 0 67896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_2_533
timestamp 1704896540
transform 1 0 73048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_2_534
timestamp 1704896540
transform 1 0 70472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_2_535
timestamp 1704896540
transform 1 0 67896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_2_536
timestamp 1704896540
transform 1 0 73048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_2_537
timestamp 1704896540
transform 1 0 70472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_2_538
timestamp 1704896540
transform 1 0 67896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_2_539
timestamp 1704896540
transform 1 0 73048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_2_540
timestamp 1704896540
transform 1 0 70472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_2_541
timestamp 1704896540
transform 1 0 67896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_2_542
timestamp 1704896540
transform 1 0 73048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_2_543
timestamp 1704896540
transform 1 0 70472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_2_544
timestamp 1704896540
transform 1 0 67896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_2_545
timestamp 1704896540
transform 1 0 73048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_2_546
timestamp 1704896540
transform 1 0 70472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_2_547
timestamp 1704896540
transform 1 0 67896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_2_548
timestamp 1704896540
transform 1 0 73048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_2_549
timestamp 1704896540
transform 1 0 70472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_2_550
timestamp 1704896540
transform 1 0 67896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_2_551
timestamp 1704896540
transform 1 0 73048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_2_552
timestamp 1704896540
transform 1 0 70472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_2_553
timestamp 1704896540
transform 1 0 67896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_2_554
timestamp 1704896540
transform 1 0 73048 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_2_555
timestamp 1704896540
transform 1 0 70472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_2_556
timestamp 1704896540
transform 1 0 67896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_2_557
timestamp 1704896540
transform 1 0 73048 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_2_558
timestamp 1704896540
transform 1 0 70472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_2_559
timestamp 1704896540
transform 1 0 67896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_2_560
timestamp 1704896540
transform 1 0 73048 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_2_561
timestamp 1704896540
transform 1 0 70472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_2_562
timestamp 1704896540
transform 1 0 67896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_2_563
timestamp 1704896540
transform 1 0 73048 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_2_564
timestamp 1704896540
transform 1 0 70472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_2_565
timestamp 1704896540
transform 1 0 67896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_2_566
timestamp 1704896540
transform 1 0 73048 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_2_567
timestamp 1704896540
transform 1 0 70472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_2_568
timestamp 1704896540
transform 1 0 67896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_2_569
timestamp 1704896540
transform 1 0 73048 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_2_570
timestamp 1704896540
transform 1 0 70472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_2_571
timestamp 1704896540
transform 1 0 67896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_2_572
timestamp 1704896540
transform 1 0 73048 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_2_573
timestamp 1704896540
transform 1 0 70472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_2_574
timestamp 1704896540
transform 1 0 67896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_2_575
timestamp 1704896540
transform 1 0 73048 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_2_576
timestamp 1704896540
transform 1 0 70472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_2_577
timestamp 1704896540
transform 1 0 67896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_2_578
timestamp 1704896540
transform 1 0 73048 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_2_579
timestamp 1704896540
transform 1 0 70472 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_2_580
timestamp 1704896540
transform 1 0 67896 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_2_581
timestamp 1704896540
transform 1 0 73048 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_2_582
timestamp 1704896540
transform 1 0 70472 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_2_583
timestamp 1704896540
transform 1 0 67896 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_2_584
timestamp 1704896540
transform 1 0 73048 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_2_585
timestamp 1704896540
transform 1 0 70472 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_2_586
timestamp 1704896540
transform 1 0 67896 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_2_587
timestamp 1704896540
transform 1 0 73048 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_2_588
timestamp 1704896540
transform 1 0 70472 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_2_589
timestamp 1704896540
transform 1 0 67896 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_2_590
timestamp 1704896540
transform 1 0 73048 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_2_591
timestamp 1704896540
transform 1 0 70472 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_2_592
timestamp 1704896540
transform 1 0 67896 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_2_593
timestamp 1704896540
transform 1 0 73048 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_2_594
timestamp 1704896540
transform 1 0 70472 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_2_595
timestamp 1704896540
transform 1 0 67896 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_2_596
timestamp 1704896540
transform 1 0 73048 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_2_597
timestamp 1704896540
transform 1 0 70472 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_2_598
timestamp 1704896540
transform 1 0 67896 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_2_599
timestamp 1704896540
transform 1 0 73048 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_2_600
timestamp 1704896540
transform 1 0 70472 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_2_601
timestamp 1704896540
transform 1 0 67896 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_2_602
timestamp 1704896540
transform 1 0 73048 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_2_603
timestamp 1704896540
transform 1 0 70472 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_2_604
timestamp 1704896540
transform 1 0 67896 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_2_605
timestamp 1704896540
transform 1 0 73048 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_103_2_606
timestamp 1704896540
transform 1 0 70472 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_2_607
timestamp 1704896540
transform 1 0 67896 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_2_608
timestamp 1704896540
transform 1 0 73048 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_105_2_609
timestamp 1704896540
transform 1 0 70472 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_2_610
timestamp 1704896540
transform 1 0 67896 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_2_611
timestamp 1704896540
transform 1 0 73048 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_2_612
timestamp 1704896540
transform 1 0 70472 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_2_613
timestamp 1704896540
transform 1 0 67896 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_2_614
timestamp 1704896540
transform 1 0 73048 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_2_615
timestamp 1704896540
transform 1 0 70472 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_2_616
timestamp 1704896540
transform 1 0 67896 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_2_617
timestamp 1704896540
transform 1 0 73048 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_2_618
timestamp 1704896540
transform 1 0 70472 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_2_619
timestamp 1704896540
transform 1 0 67896 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_2_620
timestamp 1704896540
transform 1 0 73048 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_2_621
timestamp 1704896540
transform 1 0 70472 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_2_622
timestamp 1704896540
transform 1 0 67896 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_2_623
timestamp 1704896540
transform 1 0 73048 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_2_624
timestamp 1704896540
transform 1 0 70472 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_2_625
timestamp 1704896540
transform 1 0 67896 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_2_626
timestamp 1704896540
transform 1 0 73048 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_2_627
timestamp 1704896540
transform 1 0 70472 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_2_628
timestamp 1704896540
transform 1 0 67896 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_2_629
timestamp 1704896540
transform 1 0 73048 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_2_630
timestamp 1704896540
transform 1 0 70472 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_2_631
timestamp 1704896540
transform 1 0 67896 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_2_632
timestamp 1704896540
transform 1 0 73048 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_2_633
timestamp 1704896540
transform 1 0 70472 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_2_634
timestamp 1704896540
transform 1 0 67896 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_2_635
timestamp 1704896540
transform 1 0 73048 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_2_636
timestamp 1704896540
transform 1 0 70472 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_2_637
timestamp 1704896540
transform 1 0 67896 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_2_638
timestamp 1704896540
transform 1 0 73048 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_2_639
timestamp 1704896540
transform 1 0 70472 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_2_640
timestamp 1704896540
transform 1 0 67896 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_2_641
timestamp 1704896540
transform 1 0 73048 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_2_642
timestamp 1704896540
transform 1 0 70472 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_2_643
timestamp 1704896540
transform 1 0 67896 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_2_644
timestamp 1704896540
transform 1 0 73048 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_2_645
timestamp 1704896540
transform 1 0 70472 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_2_646
timestamp 1704896540
transform 1 0 67896 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_2_647
timestamp 1704896540
transform 1 0 73048 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_2_648
timestamp 1704896540
transform 1 0 70472 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_2_649
timestamp 1704896540
transform 1 0 67896 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_2_650
timestamp 1704896540
transform 1 0 73048 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_2_651
timestamp 1704896540
transform 1 0 70472 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_2_652
timestamp 1704896540
transform 1 0 67896 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_2_653
timestamp 1704896540
transform 1 0 73048 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_2_654
timestamp 1704896540
transform 1 0 70472 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_2_655
timestamp 1704896540
transform 1 0 67896 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_2_656
timestamp 1704896540
transform 1 0 73048 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_2_657
timestamp 1704896540
transform 1 0 70472 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_2_658
timestamp 1704896540
transform 1 0 67896 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_2_659
timestamp 1704896540
transform 1 0 73048 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_139_2_660
timestamp 1704896540
transform 1 0 70472 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_140_2_661
timestamp 1704896540
transform 1 0 67896 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_140_2_662
timestamp 1704896540
transform 1 0 73048 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_141_2_663
timestamp 1704896540
transform 1 0 70472 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_142_2_664
timestamp 1704896540
transform 1 0 67896 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_142_2_665
timestamp 1704896540
transform 1 0 73048 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_143_2_666
timestamp 1704896540
transform 1 0 70472 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_144_2_667
timestamp 1704896540
transform 1 0 67896 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_144_2_668
timestamp 1704896540
transform 1 0 73048 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_145_2_669
timestamp 1704896540
transform 1 0 70472 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_2_670
timestamp 1704896540
transform 1 0 67896 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_2_671
timestamp 1704896540
transform 1 0 73048 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_2_672
timestamp 1704896540
transform 1 0 70472 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_2_673
timestamp 1704896540
transform 1 0 67896 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_2_674
timestamp 1704896540
transform 1 0 73048 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_2_675
timestamp 1704896540
transform 1 0 70472 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_2_676
timestamp 1704896540
transform 1 0 67896 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_2_677
timestamp 1704896540
transform 1 0 73048 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_2_678
timestamp 1704896540
transform 1 0 70472 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_2_679
timestamp 1704896540
transform 1 0 67896 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_2_680
timestamp 1704896540
transform 1 0 73048 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_153_2_681
timestamp 1704896540
transform 1 0 70472 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_2_682
timestamp 1704896540
transform 1 0 67896 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_2_683
timestamp 1704896540
transform 1 0 73048 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_155_2_684
timestamp 1704896540
transform 1 0 67896 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_155_2_685
timestamp 1704896540
transform 1 0 70472 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_155_2_686
timestamp 1704896540
transform 1 0 73048 0 -1 85952
box -38 -48 130 592
<< labels >>
flabel metal2 s 4188 1040 4540 5972 0 FreeSans 1792 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal2 s 14188 1040 14540 5972 0 FreeSans 1792 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal2 s 24188 1040 24540 5972 0 FreeSans 1792 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal2 s 34188 1040 34540 5972 0 FreeSans 1792 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal2 s 44188 1040 44540 5972 0 FreeSans 1792 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal2 s 54188 1040 54540 5944 0 FreeSans 1792 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal2 s 64188 1040 64540 5972 0 FreeSans 1792 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal2 s 74188 1040 74540 86000 0 FreeSans 1792 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal3 s 964 4264 75028 4616 0 FreeSans 1920 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal3 s 964 14264 75028 14616 0 FreeSans 1920 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal3 s 964 24264 75028 24616 0 FreeSans 1920 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal3 s 964 34264 75028 34616 0 FreeSans 1920 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal3 s 964 44264 75028 44616 0 FreeSans 1920 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal3 s 964 54264 75028 54616 0 FreeSans 1920 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal3 s 964 64264 75028 64616 0 FreeSans 1920 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal3 s 964 74264 75028 74616 0 FreeSans 1920 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal3 s 964 84264 75028 84616 0 FreeSans 1920 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal2 s 1836 1040 2188 5944 0 FreeSans 1792 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 11836 1040 12188 5972 0 FreeSans 1792 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 21836 1040 22188 5972 0 FreeSans 1792 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 31836 1040 32188 5972 0 FreeSans 1792 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 41836 1040 42188 5972 0 FreeSans 1792 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 51836 1040 52188 5972 0 FreeSans 1792 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 61836 1040 62188 5972 0 FreeSans 1792 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 71836 1040 72188 86000 0 FreeSans 1792 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 964 1912 75028 2264 0 FreeSans 1920 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 964 11912 75028 12264 0 FreeSans 1920 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 964 21912 75028 22264 0 FreeSans 1920 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 964 31912 75028 32264 0 FreeSans 1920 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 964 41912 75028 42264 0 FreeSans 1920 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 964 51912 75028 52264 0 FreeSans 1920 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 964 61912 75028 62264 0 FreeSans 1920 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 964 71912 75028 72264 0 FreeSans 1920 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 964 81912 75028 82264 0 FreeSans 1920 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 23018 0 23074 800 0 FreeSans 224 90 0 0 wb_clk_i
port 2 nsew signal input
flabel metal2 s 23478 0 23534 800 0 FreeSans 224 90 0 0 wb_rst_i
port 3 nsew signal input
flabel metal2 s 23938 0 23994 800 0 FreeSans 224 90 0 0 wbs_ack_o
port 4 nsew signal output
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 wbs_adr_i[0]
port 5 nsew signal input
flabel metal2 s 41418 0 41474 800 0 FreeSans 224 90 0 0 wbs_adr_i[10]
port 6 nsew signal input
flabel metal2 s 42798 0 42854 800 0 FreeSans 224 90 0 0 wbs_adr_i[11]
port 7 nsew signal input
flabel metal2 s 44178 0 44234 800 0 FreeSans 224 90 0 0 wbs_adr_i[12]
port 8 nsew signal input
flabel metal2 s 45558 0 45614 800 0 FreeSans 224 90 0 0 wbs_adr_i[13]
port 9 nsew signal input
flabel metal2 s 46938 0 46994 800 0 FreeSans 224 90 0 0 wbs_adr_i[14]
port 10 nsew signal input
flabel metal2 s 48318 0 48374 800 0 FreeSans 224 90 0 0 wbs_adr_i[15]
port 11 nsew signal input
flabel metal2 s 49698 0 49754 800 0 FreeSans 224 90 0 0 wbs_adr_i[16]
port 12 nsew signal input
flabel metal2 s 51078 0 51134 800 0 FreeSans 224 90 0 0 wbs_adr_i[17]
port 13 nsew signal input
flabel metal2 s 52458 0 52514 800 0 FreeSans 224 90 0 0 wbs_adr_i[18]
port 14 nsew signal input
flabel metal2 s 53838 0 53894 800 0 FreeSans 224 90 0 0 wbs_adr_i[19]
port 15 nsew signal input
flabel metal2 s 27618 0 27674 800 0 FreeSans 224 90 0 0 wbs_adr_i[1]
port 16 nsew signal input
flabel metal2 s 55218 0 55274 800 0 FreeSans 224 90 0 0 wbs_adr_i[20]
port 17 nsew signal input
flabel metal2 s 56598 0 56654 800 0 FreeSans 224 90 0 0 wbs_adr_i[21]
port 18 nsew signal input
flabel metal2 s 57978 0 58034 800 0 FreeSans 224 90 0 0 wbs_adr_i[22]
port 19 nsew signal input
flabel metal2 s 59358 0 59414 800 0 FreeSans 224 90 0 0 wbs_adr_i[23]
port 20 nsew signal input
flabel metal2 s 60738 0 60794 800 0 FreeSans 224 90 0 0 wbs_adr_i[24]
port 21 nsew signal input
flabel metal2 s 62118 0 62174 800 0 FreeSans 224 90 0 0 wbs_adr_i[25]
port 22 nsew signal input
flabel metal2 s 63498 0 63554 800 0 FreeSans 224 90 0 0 wbs_adr_i[26]
port 23 nsew signal input
flabel metal2 s 64878 0 64934 800 0 FreeSans 224 90 0 0 wbs_adr_i[27]
port 24 nsew signal input
flabel metal2 s 66258 0 66314 800 0 FreeSans 224 90 0 0 wbs_adr_i[28]
port 25 nsew signal input
flabel metal2 s 67638 0 67694 800 0 FreeSans 224 90 0 0 wbs_adr_i[29]
port 26 nsew signal input
flabel metal2 s 29458 0 29514 800 0 FreeSans 224 90 0 0 wbs_adr_i[2]
port 27 nsew signal input
flabel metal2 s 69018 0 69074 800 0 FreeSans 224 90 0 0 wbs_adr_i[30]
port 28 nsew signal input
flabel metal2 s 70398 0 70454 800 0 FreeSans 224 90 0 0 wbs_adr_i[31]
port 29 nsew signal input
flabel metal2 s 31298 0 31354 800 0 FreeSans 224 90 0 0 wbs_adr_i[3]
port 30 nsew signal input
flabel metal2 s 33138 0 33194 800 0 FreeSans 224 90 0 0 wbs_adr_i[4]
port 31 nsew signal input
flabel metal2 s 34518 0 34574 800 0 FreeSans 224 90 0 0 wbs_adr_i[5]
port 32 nsew signal input
flabel metal2 s 35898 0 35954 800 0 FreeSans 224 90 0 0 wbs_adr_i[6]
port 33 nsew signal input
flabel metal2 s 37278 0 37334 800 0 FreeSans 224 90 0 0 wbs_adr_i[7]
port 34 nsew signal input
flabel metal2 s 38658 0 38714 800 0 FreeSans 224 90 0 0 wbs_adr_i[8]
port 35 nsew signal input
flabel metal2 s 40038 0 40094 800 0 FreeSans 224 90 0 0 wbs_adr_i[9]
port 36 nsew signal input
flabel metal2 s 24398 0 24454 800 0 FreeSans 224 90 0 0 wbs_cyc_i
port 37 nsew signal input
flabel metal2 s 26238 0 26294 800 0 FreeSans 224 90 0 0 wbs_dat_i[0]
port 38 nsew signal input
flabel metal2 s 41878 0 41934 800 0 FreeSans 224 90 0 0 wbs_dat_i[10]
port 39 nsew signal input
flabel metal2 s 43258 0 43314 800 0 FreeSans 224 90 0 0 wbs_dat_i[11]
port 40 nsew signal input
flabel metal2 s 44638 0 44694 800 0 FreeSans 224 90 0 0 wbs_dat_i[12]
port 41 nsew signal input
flabel metal2 s 46018 0 46074 800 0 FreeSans 224 90 0 0 wbs_dat_i[13]
port 42 nsew signal input
flabel metal2 s 47398 0 47454 800 0 FreeSans 224 90 0 0 wbs_dat_i[14]
port 43 nsew signal input
flabel metal2 s 48778 0 48834 800 0 FreeSans 224 90 0 0 wbs_dat_i[15]
port 44 nsew signal input
flabel metal2 s 50158 0 50214 800 0 FreeSans 224 90 0 0 wbs_dat_i[16]
port 45 nsew signal input
flabel metal2 s 51538 0 51594 800 0 FreeSans 224 90 0 0 wbs_dat_i[17]
port 46 nsew signal input
flabel metal2 s 52918 0 52974 800 0 FreeSans 224 90 0 0 wbs_dat_i[18]
port 47 nsew signal input
flabel metal2 s 54298 0 54354 800 0 FreeSans 224 90 0 0 wbs_dat_i[19]
port 48 nsew signal input
flabel metal2 s 28078 0 28134 800 0 FreeSans 224 90 0 0 wbs_dat_i[1]
port 49 nsew signal input
flabel metal2 s 55678 0 55734 800 0 FreeSans 224 90 0 0 wbs_dat_i[20]
port 50 nsew signal input
flabel metal2 s 57058 0 57114 800 0 FreeSans 224 90 0 0 wbs_dat_i[21]
port 51 nsew signal input
flabel metal2 s 58438 0 58494 800 0 FreeSans 224 90 0 0 wbs_dat_i[22]
port 52 nsew signal input
flabel metal2 s 59818 0 59874 800 0 FreeSans 224 90 0 0 wbs_dat_i[23]
port 53 nsew signal input
flabel metal2 s 61198 0 61254 800 0 FreeSans 224 90 0 0 wbs_dat_i[24]
port 54 nsew signal input
flabel metal2 s 62578 0 62634 800 0 FreeSans 224 90 0 0 wbs_dat_i[25]
port 55 nsew signal input
flabel metal2 s 63958 0 64014 800 0 FreeSans 224 90 0 0 wbs_dat_i[26]
port 56 nsew signal input
flabel metal2 s 65338 0 65394 800 0 FreeSans 224 90 0 0 wbs_dat_i[27]
port 57 nsew signal input
flabel metal2 s 66718 0 66774 800 0 FreeSans 224 90 0 0 wbs_dat_i[28]
port 58 nsew signal input
flabel metal2 s 68098 0 68154 800 0 FreeSans 224 90 0 0 wbs_dat_i[29]
port 59 nsew signal input
flabel metal2 s 29918 0 29974 800 0 FreeSans 224 90 0 0 wbs_dat_i[2]
port 60 nsew signal input
flabel metal2 s 69478 0 69534 800 0 FreeSans 224 90 0 0 wbs_dat_i[30]
port 61 nsew signal input
flabel metal2 s 70858 0 70914 800 0 FreeSans 224 90 0 0 wbs_dat_i[31]
port 62 nsew signal input
flabel metal2 s 31758 0 31814 800 0 FreeSans 224 90 0 0 wbs_dat_i[3]
port 63 nsew signal input
flabel metal2 s 33598 0 33654 800 0 FreeSans 224 90 0 0 wbs_dat_i[4]
port 64 nsew signal input
flabel metal2 s 34978 0 35034 800 0 FreeSans 224 90 0 0 wbs_dat_i[5]
port 65 nsew signal input
flabel metal2 s 36358 0 36414 800 0 FreeSans 224 90 0 0 wbs_dat_i[6]
port 66 nsew signal input
flabel metal2 s 37738 0 37794 800 0 FreeSans 224 90 0 0 wbs_dat_i[7]
port 67 nsew signal input
flabel metal2 s 39118 0 39174 800 0 FreeSans 224 90 0 0 wbs_dat_i[8]
port 68 nsew signal input
flabel metal2 s 40498 0 40554 800 0 FreeSans 224 90 0 0 wbs_dat_i[9]
port 69 nsew signal input
flabel metal2 s 26698 0 26754 800 0 FreeSans 224 90 0 0 wbs_dat_o[0]
port 70 nsew signal output
flabel metal2 s 42338 0 42394 800 0 FreeSans 224 90 0 0 wbs_dat_o[10]
port 71 nsew signal output
flabel metal2 s 43718 0 43774 800 0 FreeSans 224 90 0 0 wbs_dat_o[11]
port 72 nsew signal output
flabel metal2 s 45098 0 45154 800 0 FreeSans 224 90 0 0 wbs_dat_o[12]
port 73 nsew signal output
flabel metal2 s 46478 0 46534 800 0 FreeSans 224 90 0 0 wbs_dat_o[13]
port 74 nsew signal output
flabel metal2 s 47858 0 47914 800 0 FreeSans 224 90 0 0 wbs_dat_o[14]
port 75 nsew signal output
flabel metal2 s 49238 0 49294 800 0 FreeSans 224 90 0 0 wbs_dat_o[15]
port 76 nsew signal output
flabel metal2 s 50618 0 50674 800 0 FreeSans 224 90 0 0 wbs_dat_o[16]
port 77 nsew signal output
flabel metal2 s 51998 0 52054 800 0 FreeSans 224 90 0 0 wbs_dat_o[17]
port 78 nsew signal output
flabel metal2 s 53378 0 53434 800 0 FreeSans 224 90 0 0 wbs_dat_o[18]
port 79 nsew signal output
flabel metal2 s 54758 0 54814 800 0 FreeSans 224 90 0 0 wbs_dat_o[19]
port 80 nsew signal output
flabel metal2 s 28538 0 28594 800 0 FreeSans 224 90 0 0 wbs_dat_o[1]
port 81 nsew signal output
flabel metal2 s 56138 0 56194 800 0 FreeSans 224 90 0 0 wbs_dat_o[20]
port 82 nsew signal output
flabel metal2 s 57518 0 57574 800 0 FreeSans 224 90 0 0 wbs_dat_o[21]
port 83 nsew signal output
flabel metal2 s 58898 0 58954 800 0 FreeSans 224 90 0 0 wbs_dat_o[22]
port 84 nsew signal output
flabel metal2 s 60278 0 60334 800 0 FreeSans 224 90 0 0 wbs_dat_o[23]
port 85 nsew signal output
flabel metal2 s 61658 0 61714 800 0 FreeSans 224 90 0 0 wbs_dat_o[24]
port 86 nsew signal output
flabel metal2 s 63038 0 63094 800 0 FreeSans 224 90 0 0 wbs_dat_o[25]
port 87 nsew signal output
flabel metal2 s 64418 0 64474 800 0 FreeSans 224 90 0 0 wbs_dat_o[26]
port 88 nsew signal output
flabel metal2 s 65798 0 65854 800 0 FreeSans 224 90 0 0 wbs_dat_o[27]
port 89 nsew signal output
flabel metal2 s 67178 0 67234 800 0 FreeSans 224 90 0 0 wbs_dat_o[28]
port 90 nsew signal output
flabel metal2 s 68558 0 68614 800 0 FreeSans 224 90 0 0 wbs_dat_o[29]
port 91 nsew signal output
flabel metal2 s 30378 0 30434 800 0 FreeSans 224 90 0 0 wbs_dat_o[2]
port 92 nsew signal output
flabel metal2 s 69938 0 69994 800 0 FreeSans 224 90 0 0 wbs_dat_o[30]
port 93 nsew signal output
flabel metal2 s 71318 0 71374 800 0 FreeSans 224 90 0 0 wbs_dat_o[31]
port 94 nsew signal output
flabel metal2 s 32218 0 32274 800 0 FreeSans 224 90 0 0 wbs_dat_o[3]
port 95 nsew signal output
flabel metal2 s 34058 0 34114 800 0 FreeSans 224 90 0 0 wbs_dat_o[4]
port 96 nsew signal output
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 wbs_dat_o[5]
port 97 nsew signal output
flabel metal2 s 36818 0 36874 800 0 FreeSans 224 90 0 0 wbs_dat_o[6]
port 98 nsew signal output
flabel metal2 s 38198 0 38254 800 0 FreeSans 224 90 0 0 wbs_dat_o[7]
port 99 nsew signal output
flabel metal2 s 39578 0 39634 800 0 FreeSans 224 90 0 0 wbs_dat_o[8]
port 100 nsew signal output
flabel metal2 s 40958 0 41014 800 0 FreeSans 224 90 0 0 wbs_dat_o[9]
port 101 nsew signal output
flabel metal2 s 27158 0 27214 800 0 FreeSans 224 90 0 0 wbs_sel_i[0]
port 102 nsew signal input
flabel metal2 s 28998 0 29054 800 0 FreeSans 224 90 0 0 wbs_sel_i[1]
port 103 nsew signal input
flabel metal2 s 30838 0 30894 800 0 FreeSans 224 90 0 0 wbs_sel_i[2]
port 104 nsew signal input
flabel metal2 s 32678 0 32734 800 0 FreeSans 224 90 0 0 wbs_sel_i[3]
port 105 nsew signal input
flabel metal2 s 24858 0 24914 800 0 FreeSans 224 90 0 0 wbs_stb_i
port 106 nsew signal input
flabel metal2 s 25318 0 25374 800 0 FreeSans 224 90 0 0 wbs_we_i
port 107 nsew signal input
rlabel via2 62636 84560 62636 84560 0 VGND
rlabel via2 62434 82208 62434 82208 0 VPWR
rlabel metal1 28152 2618 28152 2618 0 _00_
rlabel metal1 27324 2074 27324 2074 0 _01_
rlabel metal1 32246 4114 32246 4114 0 _02_
rlabel metal1 29440 2618 29440 2618 0 _03_
rlabel metal1 66286 28730 66286 28730 0 clknet_0_wb_clk_i
rlabel metal1 29578 2924 29578 2924 0 clknet_1_0__leaf_wb_clk_i
rlabel metal1 63250 53416 63250 53416 0 clknet_1_1__leaf_wb_clk_i
rlabel metal1 23874 1224 23874 1224 0 net1
rlabel metal1 39882 3570 39882 3570 0 net10
rlabel metal1 67712 37978 67712 37978 0 net100
rlabel metal2 22862 1564 22862 1564 0 net101
rlabel metal1 67850 31246 67850 31246 0 net102
rlabel metal1 43194 2618 43194 2618 0 net103
rlabel metal1 67758 18190 67758 18190 0 net104
rlabel metal1 50324 2482 50324 2482 0 net105
rlabel metal1 58374 5678 58374 5678 0 net106
rlabel metal2 67022 2652 67022 2652 0 net107
rlabel metal1 67482 38522 67482 38522 0 net108
rlabel metal2 21574 986 21574 986 0 net109
rlabel metal2 40342 3553 40342 3553 0 net11
rlabel metal1 67804 32878 67804 32878 0 net110
rlabel metal1 48714 2618 48714 2618 0 net111
rlabel metal2 56258 5542 56258 5542 0 net112
rlabel metal1 68126 2822 68126 2822 0 net113
rlabel metal1 65964 39610 65964 39610 0 net114
rlabel metal2 40342 2108 40342 2108 0 net115
rlabel metal1 67896 19822 67896 19822 0 net116
rlabel metal2 72726 2176 72726 2176 0 net117
rlabel metal1 66700 60078 66700 60078 0 net118
rlabel metal1 48668 1258 48668 1258 0 net119
rlabel metal1 24932 2278 24932 2278 0 net12
rlabel metal1 67206 13294 67206 13294 0 net120
rlabel metal1 71254 2618 71254 2618 0 net121
rlabel metal1 66424 61710 66424 61710 0 net122
rlabel metal1 38272 2958 38272 2958 0 net123
rlabel metal1 68080 21454 68080 21454 0 net124
rlabel metal1 36248 2482 36248 2482 0 net125
rlabel metal1 67850 23086 67850 23086 0 net126
rlabel metal1 46276 2618 46276 2618 0 net127
rlabel metal1 67022 14382 67022 14382 0 net128
rlabel metal2 74658 1836 74658 1836 0 net129
rlabel metal1 26542 3468 26542 3468 0 net13
rlabel metal1 67206 63342 67206 63342 0 net130
rlabel metal1 34224 2550 34224 2550 0 net131
rlabel metal1 68402 24718 68402 24718 0 net132
rlabel metal1 33810 3026 33810 3026 0 net133
rlabel metal1 68264 26894 68264 26894 0 net134
rlabel metal2 57270 1836 57270 1836 0 net135
rlabel metal2 66286 29648 66286 29648 0 net136
rlabel metal2 53038 3060 53038 3060 0 net137
rlabel metal1 66470 39950 66470 39950 0 net138
rlabel metal1 52256 2958 52256 2958 0 net139
rlabel metal1 42182 2822 42182 2822 0 net14
rlabel metal1 67758 26010 67758 26010 0 net140
rlabel metal1 25668 2482 25668 2482 0 net141
rlabel metal1 55246 5644 55246 5644 0 net142
rlabel metal1 57086 2482 57086 2482 0 net143
rlabel metal1 66378 29818 66378 29818 0 net144
rlabel metal2 27830 2652 27830 2652 0 net145
rlabel metal2 29026 2924 29026 2924 0 net146
rlabel metal2 38962 4862 38962 4862 0 net147
rlabel metal1 63250 24449 63250 24449 0 net148
rlabel metal1 59662 1326 59662 1326 0 net149
rlabel metal1 47196 1734 47196 1734 0 net15
rlabel metal1 66746 30906 66746 30906 0 net150
rlabel metal1 58374 3026 58374 3026 0 net151
rlabel metal1 67988 31994 67988 31994 0 net152
rlabel metal1 23552 1530 23552 1530 0 net153
rlabel metal1 24702 2516 24702 2516 0 net154
rlabel metal1 27232 2618 27232 2618 0 net155
rlabel metal2 31234 3468 31234 3468 0 net156
rlabel metal1 67160 27982 67160 27982 0 net157
rlabel metal2 62422 1564 62422 1564 0 net158
rlabel metal1 67620 32538 67620 32538 0 net159
rlabel metal2 47702 2040 47702 2040 0 net16
rlabel metal1 61686 2074 61686 2074 0 net160
rlabel metal1 67390 34170 67390 34170 0 net161
rlabel metal2 64998 1836 64998 1836 0 net162
rlabel metal1 67988 35258 67988 35258 0 net163
rlabel metal1 65688 3026 65688 3026 0 net164
rlabel metal1 66332 53006 66332 53006 0 net165
rlabel metal2 22678 952 22678 952 0 net166
rlabel metal1 66746 21998 66746 21998 0 net167
rlabel metal1 25254 3094 25254 3094 0 net168
rlabel metal1 27140 1938 27140 1938 0 net169
rlabel metal2 51382 4114 51382 4114 0 net17
rlabel metal2 41630 5576 41630 5576 0 net170
rlabel metal1 63250 37517 63250 37517 0 net171
rlabel metal1 23644 2618 23644 2618 0 net172
rlabel metal1 22126 1326 22126 1326 0 net173
rlabel metal1 25622 3502 25622 3502 0 net174
rlabel metal1 27830 2958 27830 2958 0 net175
rlabel metal1 66700 40494 66700 40494 0 net176
rlabel metal1 28520 1326 28520 1326 0 net177
rlabel metal1 31694 1326 31694 1326 0 net178
rlabel via2 40434 5797 40434 5797 0 net179
rlabel metal1 49496 2618 49496 2618 0 net18
rlabel metal1 63250 64446 63250 64446 0 net180
rlabel metal1 29072 1734 29072 1734 0 net181
rlabel metal2 27186 2142 27186 2142 0 net182
rlabel metal2 31326 4964 31326 4964 0 net183
rlabel metal1 32062 2482 32062 2482 0 net184
rlabel metal1 68126 35734 68126 35734 0 net185
rlabel metal1 31050 2482 31050 2482 0 net186
rlabel metal2 32982 2346 32982 2346 0 net187
rlabel metal1 64906 35666 64906 35666 0 net188
rlabel metal1 63250 81904 63250 81904 0 net189
rlabel metal2 49450 3876 49450 3876 0 net19
rlabel metal1 32476 3706 32476 3706 0 net190
rlabel metal1 32108 2550 32108 2550 0 net191
rlabel metal1 32292 2618 32292 2618 0 net192
rlabel metal1 45540 2958 45540 2958 0 net193
rlabel metal1 66700 23222 66700 23222 0 net194
rlabel metal1 43056 3366 43056 3366 0 net195
rlabel metal1 65688 22746 65688 22746 0 net196
rlabel metal1 41630 1938 41630 1938 0 net197
rlabel metal1 67436 23834 67436 23834 0 net198
rlabel metal2 39606 2108 39606 2108 0 net199
rlabel metal1 45862 2346 45862 2346 0 net2
rlabel metal1 51658 1972 51658 1972 0 net20
rlabel metal1 66608 23834 66608 23834 0 net200
rlabel metal2 36294 2210 36294 2210 0 net201
rlabel metal1 67712 24378 67712 24378 0 net202
rlabel metal2 33810 2924 33810 2924 0 net203
rlabel metal1 66562 23018 66562 23018 0 net204
rlabel metal2 36846 3468 36846 3468 0 net205
rlabel metal2 65642 24344 65642 24344 0 net206
rlabel metal1 31740 3094 31740 3094 0 net207
rlabel metal1 66286 24378 66286 24378 0 net208
rlabel metal1 29394 4114 29394 4114 0 net209
rlabel metal1 52394 3162 52394 3162 0 net21
rlabel metal1 66562 25466 66562 25466 0 net210
rlabel metal1 30406 4114 30406 4114 0 net211
rlabel metal1 66516 24650 66516 24650 0 net212
rlabel metal1 24426 3026 24426 3026 0 net213
rlabel metal1 32200 2822 32200 2822 0 net214
rlabel metal1 67436 26554 67436 26554 0 net215
rlabel metal2 20838 1054 20838 1054 0 net216
rlabel metal1 26105 2890 26105 2890 0 net217
rlabel metal2 33810 4964 33810 4964 0 net218
rlabel metal1 67712 27370 67712 27370 0 net219
rlabel metal1 59823 2618 59823 2618 0 net22
rlabel metal1 23828 3162 23828 3162 0 net220
rlabel metal1 29348 5678 29348 5678 0 net221
rlabel metal2 28474 3162 28474 3162 0 net222
rlabel metal1 29256 3094 29256 3094 0 net223
rlabel metal1 22448 1938 22448 1938 0 net224
rlabel metal2 25622 1598 25622 1598 0 net225
rlabel metal1 50784 2618 50784 2618 0 net226
rlabel metal2 51566 3026 51566 3026 0 net227
rlabel metal1 54648 4114 54648 4114 0 net228
rlabel metal1 61180 5746 61180 5746 0 net229
rlabel metal1 56258 2074 56258 2074 0 net23
rlabel metal2 48990 3332 48990 3332 0 net230
rlabel metal1 49864 2414 49864 2414 0 net231
rlabel metal1 54280 4454 54280 4454 0 net232
rlabel metal1 63250 12563 63250 12563 0 net233
rlabel metal1 49956 1938 49956 1938 0 net234
rlabel metal1 47656 3026 47656 3026 0 net235
rlabel metal1 55706 5236 55706 5236 0 net236
rlabel metal1 63250 14523 63250 14523 0 net237
rlabel metal1 47840 2414 47840 2414 0 net238
rlabel metal1 47288 1938 47288 1938 0 net239
rlabel metal2 37214 4828 37214 4828 0 net24
rlabel via2 54878 5117 54878 5117 0 net240
rlabel metal1 63250 16735 63250 16735 0 net241
rlabel metal1 45632 2618 45632 2618 0 net242
rlabel metal1 46782 2958 46782 2958 0 net243
rlabel metal2 53498 5236 53498 5236 0 net244
rlabel metal1 63250 18879 63250 18879 0 net245
rlabel metal2 43838 3468 43838 3468 0 net246
rlabel metal1 42090 2958 42090 2958 0 net247
rlabel via1 53314 4131 53314 4131 0 net248
rlabel metal1 63250 21057 63250 21057 0 net249
rlabel metal1 68632 15470 68632 15470 0 net25
rlabel metal1 42596 1530 42596 1530 0 net250
rlabel metal2 42366 3298 42366 3298 0 net251
rlabel metal2 51750 4794 51750 4794 0 net252
rlabel metal1 63250 23201 63250 23201 0 net253
rlabel metal1 39606 1190 39606 1190 0 net254
rlabel metal1 39836 2074 39836 2074 0 net255
rlabel metal2 51566 4828 51566 4828 0 net256
rlabel metal1 63250 25413 63250 25413 0 net257
rlabel metal1 36984 1938 36984 1938 0 net258
rlabel metal2 38042 3842 38042 3842 0 net259
rlabel metal1 69414 16626 69414 16626 0 net26
rlabel metal1 47886 3910 47886 3910 0 net260
rlabel metal1 63250 27693 63250 27693 0 net261
rlabel metal1 37168 3502 37168 3502 0 net262
rlabel metal2 36938 3570 36938 3570 0 net263
rlabel metal2 49358 4369 49358 4369 0 net264
rlabel metal1 63250 29735 63250 29735 0 net265
rlabel metal1 32522 1326 32522 1326 0 net266
rlabel metal1 35328 3706 35328 3706 0 net267
rlabel metal1 46046 4794 46046 4794 0 net268
rlabel metal1 63250 32015 63250 32015 0 net269
rlabel metal1 60260 2550 60260 2550 0 net27
rlabel metal1 54096 2958 54096 2958 0 net270
rlabel metal2 56718 1870 56718 1870 0 net271
rlabel metal1 67620 15130 67620 15130 0 net272
rlabel metal1 63250 54838 63250 54838 0 net273
rlabel metal2 33258 3468 33258 3468 0 net274
rlabel metal1 32890 3094 32890 3094 0 net275
rlabel metal1 42458 4454 42458 4454 0 net276
rlabel metal1 63250 34125 63250 34125 0 net277
rlabel metal1 54188 2482 54188 2482 0 net278
rlabel metal1 52348 3094 52348 3094 0 net279
rlabel metal1 68172 17646 68172 17646 0 net28
rlabel metal1 65596 27506 65596 27506 0 net280
rlabel metal1 63250 52660 63250 52660 0 net281
rlabel metal2 58466 2244 58466 2244 0 net282
rlabel metal1 58374 3094 58374 3094 0 net283
rlabel metal1 67666 15674 67666 15674 0 net284
rlabel metal1 63250 59194 63250 59194 0 net285
rlabel metal1 51888 2414 51888 2414 0 net286
rlabel metal2 51198 2414 51198 2414 0 net287
rlabel metal1 68908 25806 68908 25806 0 net288
rlabel metal1 65458 39066 65458 39066 0 net289
rlabel metal1 69092 18734 69092 18734 0 net29
rlabel metal1 55936 3502 55936 3502 0 net290
rlabel metal2 56074 2108 56074 2108 0 net291
rlabel metal1 65918 16218 65918 16218 0 net292
rlabel metal1 63250 57016 63250 57016 0 net293
rlabel metal2 61226 2108 61226 2108 0 net294
rlabel metal1 61778 1462 61778 1462 0 net295
rlabel metal1 68310 17306 68310 17306 0 net296
rlabel metal1 63250 63584 63250 63584 0 net297
rlabel metal1 29992 5134 29992 5134 0 net298
rlabel metal2 30406 4862 30406 4862 0 net299
rlabel metal1 45310 3434 45310 3434 0 net3
rlabel metal1 68126 1530 68126 1530 0 net30
rlabel via2 46690 5117 46690 5117 0 net300
rlabel metal1 63250 38699 63250 38699 0 net301
rlabel metal1 60306 1870 60306 1870 0 net302
rlabel metal2 59202 3230 59202 3230 0 net303
rlabel metal1 66746 16558 66746 16558 0 net304
rlabel metal1 63250 61372 63250 61372 0 net305
rlabel metal1 30176 2414 30176 2414 0 net306
rlabel metal1 32062 3162 32062 3162 0 net307
rlabel metal2 40618 4777 40618 4777 0 net308
rlabel metal1 63250 36303 63250 36303 0 net309
rlabel metal1 67022 20332 67022 20332 0 net31
rlabel metal2 62514 2108 62514 2108 0 net310
rlabel metal2 60766 3298 60766 3298 0 net311
rlabel metal1 67574 17850 67574 17850 0 net312
rlabel metal1 63250 65728 63250 65728 0 net313
rlabel metal1 62376 2890 62376 2890 0 net314
rlabel metal1 63940 1326 63940 1326 0 net315
rlabel metal1 67390 18938 67390 18938 0 net316
rlabel metal1 63250 67906 63250 67906 0 net317
rlabel metal1 65412 2618 65412 2618 0 net318
rlabel metal1 64584 2550 64584 2550 0 net319
rlabel metal1 68356 2006 68356 2006 0 net32
rlabel metal1 67850 20230 67850 20230 0 net320
rlabel metal1 63250 72262 63250 72262 0 net321
rlabel metal2 23506 2108 23506 2108 0 net322
rlabel metal2 23414 1088 23414 1088 0 net323
rlabel metal2 45494 5372 45494 5372 0 net324
rlabel metal1 63250 40693 63250 40693 0 net325
rlabel metal1 63848 2958 63848 2958 0 net326
rlabel metal2 67482 1530 67482 1530 0 net327
rlabel metal1 67252 19482 67252 19482 0 net328
rlabel metal1 63250 70084 63250 70084 0 net329
rlabel metal1 68080 20366 68080 20366 0 net33
rlabel metal1 66332 2958 66332 2958 0 net330
rlabel metal2 68126 2108 68126 2108 0 net331
rlabel metal1 67942 20502 67942 20502 0 net332
rlabel metal1 63250 74590 63250 74590 0 net333
rlabel metal2 21022 2108 21022 2108 0 net334
rlabel metal1 25116 3502 25116 3502 0 net335
rlabel metal2 44758 5474 44758 5474 0 net336
rlabel metal1 65918 33082 65918 33082 0 net337
rlabel metal1 69506 1326 69506 1326 0 net338
rlabel metal1 68862 3026 68862 3026 0 net339
rlabel metal1 69506 20910 69506 20910 0 net34
rlabel metal1 67344 20570 67344 20570 0 net340
rlabel metal1 63250 76618 63250 76618 0 net341
rlabel metal1 69598 2074 69598 2074 0 net342
rlabel metal1 72220 1326 72220 1326 0 net343
rlabel metal1 67988 40494 67988 40494 0 net344
rlabel metal1 63250 78796 63250 78796 0 net345
rlabel metal1 71668 2414 71668 2414 0 net346
rlabel metal2 70886 2380 70886 2380 0 net347
rlabel metal1 68632 22066 68632 22066 0 net348
rlabel metal1 63250 81008 63250 81008 0 net349
rlabel metal1 36662 5576 36662 5576 0 net35
rlabel metal2 72266 2652 72266 2652 0 net350
rlabel metal1 73876 1530 73876 1530 0 net351
rlabel metal1 69414 42670 69414 42670 0 net352
rlabel metal1 63250 83186 63250 83186 0 net353
rlabel metal1 44804 2618 44804 2618 0 net354
rlabel metal1 44988 3162 44988 3162 0 net355
rlabel metal1 55890 6800 55890 6800 0 net356
rlabel metal3 65895 41004 65895 41004 0 net357
rlabel metal1 41768 3570 41768 3570 0 net358
rlabel metal1 44160 2414 44160 2414 0 net359
rlabel metal2 71162 3774 71162 3774 0 net36
rlabel metal1 66516 22542 66516 22542 0 net360
rlabel metal1 65274 36754 65274 36754 0 net361
rlabel metal1 40756 2618 40756 2618 0 net362
rlabel metal1 40940 2074 40940 2074 0 net363
rlabel metal1 68356 23630 68356 23630 0 net364
rlabel metal1 66976 34714 66976 34714 0 net365
rlabel metal2 38778 2652 38778 2652 0 net366
rlabel metal1 39100 2074 39100 2074 0 net367
rlabel metal1 66884 23630 66884 23630 0 net368
rlabel metal1 66838 34646 66838 34646 0 net369
rlabel metal2 73462 3774 73462 3774 0 net37
rlabel metal2 35742 2108 35742 2108 0 net370
rlabel metal1 38134 2482 38134 2482 0 net371
rlabel metal1 44804 4590 44804 4590 0 net372
rlabel metal1 67068 35802 67068 35802 0 net373
rlabel metal1 34224 3570 34224 3570 0 net374
rlabel metal1 34546 2618 34546 2618 0 net375
rlabel metal1 66838 23154 66838 23154 0 net376
rlabel metal1 65872 40358 65872 40358 0 net377
rlabel metal2 36018 3604 36018 3604 0 net378
rlabel metal1 36340 3162 36340 3162 0 net379
rlabel metal2 39974 4828 39974 4828 0 net38
rlabel metal2 66608 20060 66608 20060 0 net380
rlabel metal1 65366 34714 65366 34714 0 net381
rlabel metal1 30314 2618 30314 2618 0 net382
rlabel metal1 30038 3536 30038 3536 0 net383
rlabel metal2 66516 20332 66516 20332 0 net384
rlabel metal1 65596 36890 65596 36890 0 net385
rlabel metal1 29578 3706 29578 3706 0 net386
rlabel metal2 29670 4318 29670 4318 0 net387
rlabel via2 39514 5899 39514 5899 0 net388
rlabel metal1 65274 36346 65274 36346 0 net389
rlabel metal2 40250 3842 40250 3842 0 net39
rlabel metal2 28658 3434 28658 3434 0 net390
rlabel metal1 29072 4114 29072 4114 0 net391
rlabel via2 38778 5661 38778 5661 0 net392
rlabel metal1 65320 44710 65320 44710 0 net393
rlabel metal1 22908 2618 22908 2618 0 net394
rlabel metal2 26726 3162 26726 3162 0 net395
rlabel metal1 29762 3094 29762 3094 0 net396
rlabel metal1 20286 1292 20286 1292 0 net397
rlabel metal1 24334 2448 24334 2448 0 net398
rlabel metal1 32936 4114 32936 4114 0 net399
rlabel metal2 38134 5474 38134 5474 0 net4
rlabel metal1 42274 4726 42274 4726 0 net40
rlabel metal2 36478 5508 36478 5508 0 net400
rlabel metal2 27370 4012 27370 4012 0 net401
rlabel metal1 23552 2006 23552 2006 0 net402
rlabel metal1 21988 2074 21988 2074 0 net403
rlabel metal1 25530 1938 25530 1938 0 net404
rlabel metal2 51382 2652 51382 2652 0 net405
rlabel metal2 50462 3196 50462 3196 0 net406
rlabel metal1 51566 1360 51566 1360 0 net407
rlabel metal1 48300 3502 48300 3502 0 net408
rlabel metal2 47518 3332 47518 3332 0 net409
rlabel metal2 36754 4352 36754 4352 0 net41
rlabel metal2 49450 2210 49450 2210 0 net410
rlabel metal1 46736 3434 46736 3434 0 net411
rlabel metal1 49036 1394 49036 1394 0 net412
rlabel metal2 46138 2244 46138 2244 0 net413
rlabel metal1 46276 3366 46276 3366 0 net414
rlabel metal1 43424 3706 43424 3706 0 net415
rlabel metal1 45218 2822 45218 2822 0 net416
rlabel metal1 44666 1326 44666 1326 0 net417
rlabel metal1 42642 2482 42642 2482 0 net418
rlabel metal1 38272 1326 38272 1326 0 net419
rlabel metal2 37950 4318 37950 4318 0 net42
rlabel metal1 40480 2414 40480 2414 0 net420
rlabel metal1 38042 2618 38042 2618 0 net421
rlabel metal1 37168 2074 37168 2074 0 net422
rlabel metal2 36110 3060 36110 3060 0 net423
rlabel metal2 35650 3230 35650 3230 0 net424
rlabel metal1 34868 3162 34868 3162 0 net425
rlabel metal1 32890 1530 32890 1530 0 net426
rlabel metal1 54234 3026 54234 3026 0 net427
rlabel metal1 55016 2822 55016 2822 0 net428
rlabel metal1 30452 1190 30452 1190 0 net429
rlabel metal1 42274 3128 42274 3128 0 net43
rlabel metal2 32614 3332 32614 3332 0 net430
rlabel metal2 52670 3332 52670 3332 0 net431
rlabel metal1 53728 2414 53728 2414 0 net432
rlabel metal1 56074 2890 56074 2890 0 net433
rlabel metal2 55614 3196 55614 3196 0 net434
rlabel metal1 57408 1870 57408 1870 0 net435
rlabel metal1 57868 2414 57868 2414 0 net436
rlabel metal1 54050 1190 54050 1190 0 net437
rlabel metal2 53222 2108 53222 2108 0 net438
rlabel metal1 58696 2822 58696 2822 0 net439
rlabel metal2 40894 3689 40894 3689 0 net44
rlabel metal1 60444 2074 60444 2074 0 net440
rlabel metal1 60168 2482 60168 2482 0 net441
rlabel metal1 29440 2482 29440 2482 0 net442
rlabel metal1 60904 2822 60904 2822 0 net443
rlabel metal2 29394 5372 29394 5372 0 net444
rlabel metal1 61732 2550 61732 2550 0 net445
rlabel metal1 63296 2958 63296 2958 0 net446
rlabel metal1 24150 2380 24150 2380 0 net447
rlabel metal2 66102 2244 66102 2244 0 net448
rlabel metal2 26174 4964 26174 4964 0 net449
rlabel metal2 36570 3570 36570 3570 0 net45
rlabel metal1 66010 2822 66010 2822 0 net450
rlabel metal1 69966 1326 69966 1326 0 net451
rlabel metal2 70702 2108 70702 2108 0 net452
rlabel metal2 70702 2686 70702 2686 0 net453
rlabel metal2 73278 2142 73278 2142 0 net454
rlabel metal1 46138 1530 46138 1530 0 net455
rlabel metal1 42504 3706 42504 3706 0 net456
rlabel metal1 41676 2482 41676 2482 0 net457
rlabel metal1 40710 1258 40710 1258 0 net458
rlabel metal1 35512 1530 35512 1530 0 net459
rlabel metal1 37766 4080 37766 4080 0 net46
rlabel metal1 33948 2278 33948 2278 0 net460
rlabel metal2 34914 3196 34914 3196 0 net461
rlabel metal2 30774 2958 30774 2958 0 net462
rlabel metal2 25438 2618 25438 2618 0 net463
rlabel metal1 28750 3468 28750 3468 0 net464
rlabel metal2 36570 1122 36570 1122 0 net47
rlabel metal2 40434 3298 40434 3298 0 net48
rlabel metal2 26266 3332 26266 3332 0 net49
rlabel metal2 36110 4828 36110 4828 0 net5
rlabel metal2 26450 2414 26450 2414 0 net50
rlabel metal1 28934 2822 28934 2822 0 net51
rlabel metal2 63894 1836 63894 1836 0 net52
rlabel metal2 59754 1972 59754 1972 0 net53
rlabel metal1 63250 19243 63250 19243 0 net54
rlabel metal1 63441 17110 63441 17110 0 net55
rlabel metal1 63250 14921 63250 14921 0 net56
rlabel metal1 64407 12750 64407 12750 0 net57
rlabel metal2 51474 816 51474 816 0 net58
rlabel metal1 52210 1938 52210 1938 0 net59
rlabel metal2 40158 4420 40158 4420 0 net6
rlabel metal1 63250 52466 63250 52466 0 net60
rlabel metal1 56074 1836 56074 1836 0 net61
rlabel metal1 56534 1258 56534 1258 0 net62
rlabel metal1 63250 41023 63250 41023 0 net63
rlabel metal1 63250 59048 63250 59048 0 net64
rlabel metal1 63395 61204 63395 61204 0 net65
rlabel metal1 60444 1938 60444 1938 0 net66
rlabel metal1 62054 1326 62054 1326 0 net67
rlabel metal2 63158 850 63158 850 0 net68
rlabel metal1 63756 1938 63756 1938 0 net69
rlabel metal1 36478 4556 36478 4556 0 net7
rlabel metal1 63250 71932 63250 71932 0 net70
rlabel metal1 63250 74178 63250 74178 0 net71
rlabel metal1 63250 76472 63250 76472 0 net72
rlabel metal1 63250 78636 63250 78636 0 net73
rlabel metal1 63349 38910 63349 38910 0 net74
rlabel metal1 63250 80814 63250 80814 0 net75
rlabel metal1 63250 82992 63250 82992 0 net76
rlabel metal1 63250 36633 63250 36633 0 net77
rlabel metal1 60030 1496 60030 1496 0 net78
rlabel metal2 36938 986 36938 986 0 net79
rlabel metal1 37030 4658 37030 4658 0 net8
rlabel metal1 38594 1972 38594 1972 0 net80
rlabel metal2 39422 952 39422 952 0 net81
rlabel metal2 41170 1156 41170 1156 0 net82
rlabel metal1 63250 23565 63250 23565 0 net83
rlabel metal1 63158 49590 63158 49590 0 net84
rlabel metal1 63250 43679 63250 43679 0 net85
rlabel metal1 63250 42543 63250 42543 0 net86
rlabel metal1 63250 50114 63250 50114 0 net87
rlabel metal1 63441 52094 63441 52094 0 net88
rlabel metal1 63250 52289 63250 52289 0 net89
rlabel metal1 37674 4012 37674 4012 0 net9
rlabel metal1 63349 48715 63349 48715 0 net90
rlabel metal1 69184 15334 69184 15334 0 net91
rlabel metal2 70886 27642 70886 27642 0 net92
rlabel metal1 51612 2482 51612 2482 0 net93
rlabel metal1 58696 5338 58696 5338 0 net94
rlabel metal1 30820 4114 30820 4114 0 net95
rlabel metal1 66746 30158 66746 30158 0 net96
rlabel metal1 44574 2890 44574 2890 0 net97
rlabel metal1 66010 15334 66010 15334 0 net98
rlabel metal1 64814 2822 64814 2822 0 net99
rlabel metal2 36754 6086 36754 6086 0 ram_controller.EN
rlabel metal1 40526 4692 40526 4692 0 ram_controller.R_WB
rlabel metal2 23046 2047 23046 2047 0 wb_clk_i
rlabel metal2 23506 823 23506 823 0 wb_rst_i
rlabel metal2 23966 1010 23966 1010 0 wbs_ack_o
rlabel metal2 41446 1095 41446 1095 0 wbs_adr_i[10]
rlabel metal2 42826 1078 42826 1078 0 wbs_adr_i[11]
rlabel metal2 29486 1112 29486 1112 0 wbs_adr_i[2]
rlabel metal2 31326 2676 31326 2676 0 wbs_adr_i[3]
rlabel metal2 33166 2098 33166 2098 0 wbs_adr_i[4]
rlabel metal2 34546 823 34546 823 0 wbs_adr_i[5]
rlabel metal2 35926 2132 35926 2132 0 wbs_adr_i[6]
rlabel metal2 37306 1010 37306 1010 0 wbs_adr_i[7]
rlabel metal2 38686 1078 38686 1078 0 wbs_adr_i[8]
rlabel metal2 40066 1894 40066 1894 0 wbs_adr_i[9]
rlabel metal2 24426 823 24426 823 0 wbs_cyc_i
rlabel metal2 26266 1367 26266 1367 0 wbs_dat_i[0]
rlabel metal2 41906 823 41906 823 0 wbs_dat_i[10]
rlabel metal2 43286 1248 43286 1248 0 wbs_dat_i[11]
rlabel metal2 44666 1095 44666 1095 0 wbs_dat_i[12]
rlabel metal1 47058 2890 47058 2890 0 wbs_dat_i[13]
rlabel metal1 51888 1326 51888 1326 0 wbs_dat_i[14]
rlabel metal2 48806 1027 48806 1027 0 wbs_dat_i[15]
rlabel metal1 51658 1224 51658 1224 0 wbs_dat_i[16]
rlabel metal2 51566 959 51566 959 0 wbs_dat_i[17]
rlabel metal1 55430 1938 55430 1938 0 wbs_dat_i[18]
rlabel metal2 54326 823 54326 823 0 wbs_dat_i[19]
rlabel metal1 25737 3026 25737 3026 0 wbs_dat_i[1]
rlabel metal1 56028 2958 56028 2958 0 wbs_dat_i[20]
rlabel metal1 57454 2958 57454 2958 0 wbs_dat_i[21]
rlabel metal2 58466 1146 58466 1146 0 wbs_dat_i[22]
rlabel metal1 59938 2958 59938 2958 0 wbs_dat_i[23]
rlabel metal2 61226 823 61226 823 0 wbs_dat_i[24]
rlabel metal2 62606 1010 62606 1010 0 wbs_dat_i[25]
rlabel metal2 63986 1282 63986 1282 0 wbs_dat_i[26]
rlabel metal2 65366 1588 65366 1588 0 wbs_dat_i[27]
rlabel metal2 66746 823 66746 823 0 wbs_dat_i[28]
rlabel metal2 68126 823 68126 823 0 wbs_dat_i[29]
rlabel metal2 29946 2234 29946 2234 0 wbs_dat_i[2]
rlabel metal1 69598 2958 69598 2958 0 wbs_dat_i[30]
rlabel metal2 70886 1010 70886 1010 0 wbs_dat_i[31]
rlabel metal2 31786 2115 31786 2115 0 wbs_dat_i[3]
rlabel metal2 33626 806 33626 806 0 wbs_dat_i[4]
rlabel metal2 35006 1860 35006 1860 0 wbs_dat_i[5]
rlabel metal2 36386 1588 36386 1588 0 wbs_dat_i[6]
rlabel metal2 37766 1588 37766 1588 0 wbs_dat_i[7]
rlabel metal2 39146 1316 39146 1316 0 wbs_dat_i[8]
rlabel metal2 40526 823 40526 823 0 wbs_dat_i[9]
rlabel metal2 26726 959 26726 959 0 wbs_dat_o[0]
rlabel metal2 42366 1316 42366 1316 0 wbs_dat_o[10]
rlabel metal2 43746 1316 43746 1316 0 wbs_dat_o[11]
rlabel metal2 45126 1010 45126 1010 0 wbs_dat_o[12]
rlabel metal2 46506 1010 46506 1010 0 wbs_dat_o[13]
rlabel metal2 47886 1316 47886 1316 0 wbs_dat_o[14]
rlabel metal2 49266 1010 49266 1010 0 wbs_dat_o[15]
rlabel metal2 50646 1316 50646 1316 0 wbs_dat_o[16]
rlabel metal2 52026 823 52026 823 0 wbs_dat_o[17]
rlabel metal2 53406 1316 53406 1316 0 wbs_dat_o[18]
rlabel metal2 54786 1010 54786 1010 0 wbs_dat_o[19]
rlabel metal2 28566 1010 28566 1010 0 wbs_dat_o[1]
rlabel metal2 56166 1316 56166 1316 0 wbs_dat_o[20]
rlabel metal2 57546 1010 57546 1010 0 wbs_dat_o[21]
rlabel metal2 58926 1316 58926 1316 0 wbs_dat_o[22]
rlabel metal2 60306 1010 60306 1010 0 wbs_dat_o[23]
rlabel metal2 61686 1010 61686 1010 0 wbs_dat_o[24]
rlabel metal2 63066 1316 63066 1316 0 wbs_dat_o[25]
rlabel metal2 64446 823 64446 823 0 wbs_dat_o[26]
rlabel metal2 65826 1010 65826 1010 0 wbs_dat_o[27]
rlabel metal2 67206 1078 67206 1078 0 wbs_dat_o[28]
rlabel metal2 68586 1316 68586 1316 0 wbs_dat_o[29]
rlabel metal2 30406 1316 30406 1316 0 wbs_dat_o[2]
rlabel metal2 69966 1078 69966 1078 0 wbs_dat_o[30]
rlabel metal2 71346 1316 71346 1316 0 wbs_dat_o[31]
rlabel metal2 32246 1316 32246 1316 0 wbs_dat_o[3]
rlabel metal2 34086 1316 34086 1316 0 wbs_dat_o[4]
rlabel metal2 35466 1010 35466 1010 0 wbs_dat_o[5]
rlabel metal2 36846 1316 36846 1316 0 wbs_dat_o[6]
rlabel metal2 38226 1010 38226 1010 0 wbs_dat_o[7]
rlabel metal2 39606 1010 39606 1010 0 wbs_dat_o[8]
rlabel metal2 40986 823 40986 823 0 wbs_dat_o[9]
rlabel metal1 25346 2380 25346 2380 0 wbs_sel_i[0]
rlabel metal2 25162 1054 25162 1054 0 wbs_sel_i[1]
rlabel metal2 26174 1666 26174 1666 0 wbs_sel_i[2]
rlabel metal2 32706 1299 32706 1299 0 wbs_sel_i[3]
rlabel metal2 24886 1248 24886 1248 0 wbs_stb_i
rlabel metal2 25346 1316 25346 1316 0 wbs_we_i
<< properties >>
string FIXED_BBOX 0 0 76000 87000
<< end >>
